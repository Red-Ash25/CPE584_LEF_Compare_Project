# 
# LEF OUT 
# User Name : iptguser 
# Date : Mon Feb  4 15:39:10 2013
# 
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO scs8ls_tapvgndnovpb_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.48 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.48 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.48 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb
  OBS
    LAYER li1 ;
      RECT 0 3.245 0.48 3.415 ;
      RECT 0.09 0.085 0.39 1.44 ;
      RECT 0 -0.085 0.48 0.085 ;
    LAYER mcon ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_tapvgndnovpb_1

MACRO scs8ls_decaphe_18
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 0.085 1.77 8.555 3.245 ;
      RECT 1.325 1.25 2.015 1.77 ;
      RECT 3.085 1.25 3.775 1.77 ;
      RECT 4.845 1.25 5.535 1.77 ;
      RECT 6.605 1.25 7.295 1.77 ;
      RECT 0.085 1.08 1.155 1.6 ;
      RECT 0.085 0.085 8.555 1.08 ;
      RECT 2.205 1.08 2.895 1.6 ;
      RECT 3.965 1.08 4.655 1.6 ;
      RECT 5.725 1.08 6.415 1.6 ;
      RECT 7.485 1.08 8.555 1.6 ;
      RECT 0 -0.085 8.64 0.085 ;
    LAYER mcon ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
  END
END scs8ls_decaphe_18

MACRO scs8ls_decaphe_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.96 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.96 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.96 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 0.96 3.415 ;
      RECT 0.085 1.845 0.875 3.245 ;
      RECT 0.085 0.085 0.47 1.675 ;
      RECT 0 -0.085 0.96 0.085 ;
    LAYER mcon ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_decaphe_2

MACRO scs8ls_decaphe_3
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 1.44 3.415 ;
      RECT 0.085 1.77 1.355 3.245 ;
      RECT 0.805 1.25 1.355 1.77 ;
      RECT 0.085 1.08 0.635 1.6 ;
      RECT 0.085 0.085 1.355 1.08 ;
      RECT 0 -0.085 1.44 0.085 ;
    LAYER mcon ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
  END
END scs8ls_decaphe_3

MACRO scs8ls_decaphe_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 1.92 3.415 ;
      RECT 0.085 1.77 1.835 3.245 ;
      RECT 1.06 1.25 1.835 1.77 ;
      RECT 0.085 1.08 0.89 1.6 ;
      RECT 0.085 0.085 1.835 1.08 ;
      RECT 0 -0.085 1.92 0.085 ;
    LAYER mcon ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
  END
END scs8ls_decaphe_4

MACRO scs8ls_decaphe_6
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 0.12 1.77 2.76 3.245 ;
      RECT 1.365 1.25 2.76 1.77 ;
      RECT 0.12 1.08 1.195 1.6 ;
      RECT 0.12 0.085 2.76 1.08 ;
      RECT 0 -0.085 2.88 0.085 ;
    LAYER mcon ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
  END
END scs8ls_decaphe_6

MACRO scs8ls_decaphe_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.085 1.075 0.95 1.6 ;
      RECT 0.085 1.07 2.71 1.075 ;
      RECT 2 1.075 2.71 1.6 ;
      RECT 0.085 0.085 3.755 1.07 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 0.085 1.77 3.755 3.245 ;
      RECT 1.12 1.25 1.83 1.77 ;
      RECT 2.88 1.25 3.755 1.77 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_decaphe_8

MACRO scs8ls_fill_diode_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 0.135 0.085 3.705 0.58 ;
      RECT 0.135 2.75 3.705 3.245 ;
      RECT 0 3.245 3.84 3.415 ;
    LAYER mcon ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
  END
END scs8ls_fill_diode_8

MACRO scs8ls_fill_diode_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.92 0.085 ;
      RECT 0.135 0.085 1.785 0.58 ;
      RECT 0.135 2.75 1.785 3.245 ;
      RECT 0 3.245 1.92 3.415 ;
    LAYER mcon ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
  END
END scs8ls_fill_diode_4

MACRO scs8ls_fill_diode_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.96 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.96 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 0.96 0.085 ;
      RECT 0.135 0.085 0.825 0.58 ;
      RECT 0.135 2.75 0.825 3.245 ;
      RECT 0 3.245 0.96 3.415 ;
    LAYER mcon ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_fill_diode_2

MACRO scs8ls_diode_2
  CLASS CORE ANTENNACELL ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.96 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.96 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb

  PIN DIODE
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.265 0.865 3.065 ;
    END
    ANTENNADIFFAREA 0.6417 ;
  END DIODE
  OBS
    LAYER li1 ;
      RECT 0 -0.085 0.96 0.085 ;
      RECT 0 3.245 0.96 3.415 ;
    LAYER mcon ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_diode_2

MACRO scs8ls_tapmet1_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.96 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.96 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.56 2.645 0.88 2.905 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.08 0.425 0.4 0.685 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.09 0.265 0.87 1.105 ;
      RECT 0 -0.085 0.96 0.085 ;
      RECT 0 3.245 0.96 3.415 ;
      RECT 0.09 2.21 0.87 3.065 ;
    LAYER mcon ;
      RECT 0.635 2.69 0.805 2.86 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 0.47 0.325 0.64 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_tapmet1_2

MACRO scs8ls_sedfxbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 17.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.45 1.905 1.78 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END DE

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.475 1.18 4.915 1.51 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.125 1.18 5.635 1.51 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.705 1.18 7.045 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.98 0.835 1.99 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.355 0.35 16.685 0.96 ;
        RECT 16.355 0.96 17.165 1.13 ;
        RECT 16.7 1.13 17.165 1.805 ;
        RECT 16.435 1.805 17.165 1.975 ;
        RECT 16.435 1.975 16.665 3.01 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.485 0.35 15.825 2.15 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 17.28 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 17.28 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 7.215 1.01 7.385 1.47 ;
      RECT 6.915 0.35 7.385 1.01 ;
      RECT 4.055 1.68 6.135 1.85 ;
      RECT 5.805 1.85 6.135 2.085 ;
      RECT 5.805 1.43 6.135 1.68 ;
      RECT 4.135 2.245 4.525 2.735 ;
      RECT 4.055 0.605 4.79 1.01 ;
      RECT 4.135 2.055 4.305 2.245 ;
      RECT 4.055 1.85 4.305 2.055 ;
      RECT 4.055 1.01 4.305 1.68 ;
      RECT 4.055 0.365 4.305 0.605 ;
      RECT 0.085 2.29 1.655 2.46 ;
      RECT 1.485 2.46 1.655 2.905 ;
      RECT 1.485 2.905 2.335 3.075 ;
      RECT 2.165 2.46 2.335 2.905 ;
      RECT 2.165 2.29 3.545 2.46 ;
      RECT 3.265 2.46 3.545 2.97 ;
      RECT 3.375 1.345 3.545 2.29 ;
      RECT 3 1.175 3.545 1.345 ;
      RECT 3 0.545 3.33 1.175 ;
      RECT 0.085 2.46 0.525 2.98 ;
      RECT 0.085 0.42 0.58 0.73 ;
      RECT 0.085 0.73 0.255 2.29 ;
      RECT 2.875 1.515 3.205 1.845 ;
      RECT 1.825 2.12 1.995 2.735 ;
      RECT 1.005 1.95 2.635 2.12 ;
      RECT 2.305 1.515 2.635 1.95 ;
      RECT 1.005 1.11 2.01 1.28 ;
      RECT 1.68 0.545 2.01 1.11 ;
      RECT 1.005 1.28 1.335 1.95 ;
      RECT 15.995 1.3 16.51 1.635 ;
      RECT 14.475 2.38 16.185 2.49 ;
      RECT 13.585 2.32 16.185 2.38 ;
      RECT 15.995 1.635 16.185 2.32 ;
      RECT 14.475 2.49 14.835 2.98 ;
      RECT 13.585 2.055 15.235 2.32 ;
      RECT 14.475 1.8 15.235 2.055 ;
      RECT 14.665 1.55 15.235 1.8 ;
      RECT 14.665 1.13 14.835 1.55 ;
      RECT 14.505 0.35 14.835 1.13 ;
      RECT 0 3.245 17.28 3.415 ;
      RECT 16.835 2.145 17.165 3.245 ;
      RECT 15.935 2.66 16.265 3.245 ;
      RECT 10.225 2.73 10.555 3.245 ;
      RECT 11.32 2.73 11.65 3.245 ;
      RECT 15.035 2.66 15.365 3.245 ;
      RECT 6.485 2.65 6.735 3.245 ;
      RECT 7.795 2.65 8.125 3.245 ;
      RECT 13.765 2.65 14.305 3.245 ;
      RECT 1.065 2.63 1.315 3.245 ;
      RECT 2.505 2.63 2.755 3.245 ;
      RECT 5.035 2.595 5.305 3.245 ;
      RECT 12.89 2.52 13.325 2.98 ;
      RECT 13.155 1.885 13.325 2.52 ;
      RECT 13.155 1.715 13.865 1.885 ;
      RECT 13.695 1.63 13.865 1.715 ;
      RECT 13.695 1.3 14.495 1.63 ;
      RECT 13.695 0.94 13.865 1.3 ;
      RECT 12.42 0.77 13.865 0.94 ;
      RECT 12.42 0.35 12.75 0.77 ;
      RECT 8.725 2.14 9.055 2.305 ;
      RECT 8.245 1.82 9.055 2.14 ;
      RECT 8.885 0.425 9.055 1.82 ;
      RECT 7.905 0.255 9.735 0.425 ;
      RECT 7.905 0.425 8.235 1.13 ;
      RECT 9.565 0.425 9.735 0.85 ;
      RECT 9.565 0.85 10.86 1.02 ;
      RECT 9.565 1.02 9.855 1.345 ;
      RECT 10.69 0.425 10.86 0.85 ;
      RECT 10.69 0.255 11.54 0.425 ;
      RECT 11.37 0.425 11.54 0.85 ;
      RECT 11.37 0.85 12.25 1.02 ;
      RECT 12.08 1.02 12.25 1.13 ;
      RECT 12.08 1.13 13.525 1.3 ;
      RECT 12.08 1.3 12.38 1.8 ;
      RECT 13.195 1.3 13.525 1.545 ;
      RECT 9.755 2.39 12.72 2.56 ;
      RECT 9.755 2.36 9.925 2.39 ;
      RECT 12.55 1.8 12.72 2.39 ;
      RECT 9.565 2.03 9.925 2.36 ;
      RECT 12.55 1.47 12.985 1.8 ;
      RECT 10.76 2.05 11.385 2.22 ;
      RECT 11.215 1.52 11.385 2.05 ;
      RECT 11.215 1.36 11.885 1.52 ;
      RECT 10.065 1.19 11.885 1.36 ;
      RECT 10.065 1.36 10.395 1.52 ;
      RECT 11.03 0.595 11.2 1.19 ;
      RECT 9.225 2.53 9.585 2.98 ;
      RECT 9.225 1.86 9.395 2.53 ;
      RECT 9.225 1.69 10.94 1.86 ;
      RECT 10.61 1.53 10.94 1.69 ;
      RECT 9.225 0.595 9.395 1.69 ;
      RECT 4.695 2.31 8.465 2.425 ;
      RECT 5.845 2.425 8.465 2.48 ;
      RECT 7.905 1.65 8.075 2.31 ;
      RECT 8.295 2.48 9.055 2.65 ;
      RECT 7.905 1.48 8.715 1.65 ;
      RECT 8.805 2.65 9.055 2.98 ;
      RECT 8.465 0.595 8.715 1.48 ;
      RECT 4.695 2.255 6.475 2.31 ;
      RECT 5.845 2.48 6.305 2.925 ;
      RECT 6.305 1.26 6.475 2.255 ;
      RECT 5.82 1.09 6.475 1.26 ;
      RECT 5.82 0.605 6.15 1.09 ;
      RECT 3.715 2.905 4.865 3.075 ;
      RECT 4.695 2.425 4.865 2.905 ;
      RECT 3.715 2.29 3.965 2.905 ;
      RECT 3.715 1.005 3.885 2.29 ;
      RECT 3.5 0.545 3.885 1.005 ;
      RECT 0 -0.085 17.28 0.085 ;
      RECT 16.855 0.085 17.115 0.79 ;
      RECT 16.005 0.085 16.175 1.13 ;
      RECT 14.065 0.6 14.335 1.12 ;
      RECT 13.32 0.085 14.335 0.6 ;
      RECT 1.07 0.085 1.4 0.81 ;
      RECT 2.18 0.085 2.51 1.005 ;
      RECT 4.96 0.085 5.29 1.01 ;
      RECT 6.415 0.085 6.745 0.92 ;
      RECT 7.555 0.085 7.725 1.13 ;
      RECT 10.27 0.085 10.52 0.68 ;
      RECT 11.71 0.085 11.96 0.68 ;
      RECT 15.065 0.085 15.315 1.13 ;
      RECT 6.855 1.82 7.655 2.14 ;
      RECT 7.215 1.47 7.655 1.82 ;
    LAYER mcon ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 1.58 3.205 1.75 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 16.955 -0.085 17.125 0.085 ;
      RECT 16.955 3.245 17.125 3.415 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 1.58 15.205 1.75 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
    LAYER met1 ;
      RECT 2.975 1.735 3.265 1.78 ;
      RECT 2.975 1.595 15.265 1.735 ;
      RECT 14.975 1.735 15.265 1.78 ;
      RECT 2.975 1.55 3.265 1.595 ;
      RECT 14.975 1.55 15.265 1.595 ;
  END
END scs8ls_sedfxbp_2

MACRO scs8ls_sedfxtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 15.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.11 0.805 1.78 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515 1.32 1.845 1.78 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END DE

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.4 1.18 4.73 1.51 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.18 5.28 1.745 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.475 0.35 14.815 2.98 ;
    END
    ANTENNADIFFAREA 0.5189 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.33 1.18 6.66 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 15.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 15.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 14.075 1.58 14.245 1.75 ;
      RECT 2.555 1.58 2.725 1.75 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
    LAYER met1 ;
      RECT 2.495 1.735 2.785 1.78 ;
      RECT 2.495 1.595 14.305 1.735 ;
      RECT 14.015 1.735 14.305 1.78 ;
      RECT 2.495 1.55 2.785 1.595 ;
      RECT 14.015 1.55 14.305 1.595 ;
    LAYER li1 ;
      RECT 8.985 2.56 9.315 2.98 ;
      RECT 8.835 2.39 9.315 2.56 ;
      RECT 8.835 1.79 9.005 2.39 ;
      RECT 8.745 1.62 10.465 1.79 ;
      RECT 10.135 1.79 10.465 1.795 ;
      RECT 10.135 1.535 10.465 1.62 ;
      RECT 8.745 0.595 8.915 1.62 ;
      RECT 1.705 2.12 1.875 2.735 ;
      RECT 0.975 1.95 2.385 2.12 ;
      RECT 2.055 1.52 2.385 1.95 ;
      RECT 0.975 0.995 1.81 1.15 ;
      RECT 0.975 0.98 1.89 0.995 ;
      RECT 1.64 0.535 1.89 0.98 ;
      RECT 0.975 1.15 1.305 1.95 ;
      RECT 9.485 2.39 12.2 2.56 ;
      RECT 9.485 2.22 9.655 2.39 ;
      RECT 12.03 1.735 12.2 2.39 ;
      RECT 9.175 1.96 9.655 2.22 ;
      RECT 12.03 1.45 12.465 1.735 ;
      RECT 3.905 1.915 5.82 2.085 ;
      RECT 5.49 1.415 5.82 1.915 ;
      RECT 3.905 0.605 4.575 1.01 ;
      RECT 4.015 2.255 4.37 2.735 ;
      RECT 4.015 2.085 4.185 2.255 ;
      RECT 3.905 1.01 4.185 1.915 ;
      RECT 3.905 0.255 4.185 0.605 ;
      RECT 12.37 1.94 12.805 2.98 ;
      RECT 12.635 1.905 12.805 1.94 ;
      RECT 12.635 1.735 13.785 1.905 ;
      RECT 13.615 1.38 13.785 1.735 ;
      RECT 13.175 0.94 13.345 1.735 ;
      RECT 13.615 1.05 13.945 1.38 ;
      RECT 11.9 0.77 13.345 0.94 ;
      RECT 11.9 0.35 12.23 0.77 ;
      RECT 6.61 1.83 7.39 2.16 ;
      RECT 6.61 1.76 7 1.83 ;
      RECT 6.83 1.01 7 1.76 ;
      RECT 6.45 0.84 7 1.01 ;
      RECT 6.45 0.35 6.78 0.84 ;
      RECT 2.555 1.505 3.055 1.835 ;
      RECT 10.385 1.97 10.805 2.22 ;
      RECT 10.635 1.525 10.805 1.97 ;
      RECT 10.635 1.365 11.385 1.525 ;
      RECT 9.565 1.195 11.385 1.365 ;
      RECT 9.565 1.365 9.895 1.45 ;
      RECT 9.565 1.19 9.895 1.195 ;
      RECT 10.51 0.595 10.68 1.195 ;
      RECT 0.085 2.29 1.535 2.46 ;
      RECT 1.365 2.46 1.535 2.905 ;
      RECT 1.365 2.905 2.215 3.075 ;
      RECT 2.045 2.46 2.215 2.905 ;
      RECT 2.045 2.29 3.395 2.46 ;
      RECT 3.145 2.46 3.395 2.975 ;
      RECT 3.225 1.335 3.395 2.29 ;
      RECT 2.89 1.165 3.395 1.335 ;
      RECT 2.89 0.535 3.22 1.165 ;
      RECT 0.085 2.46 0.435 2.98 ;
      RECT 0.085 0.48 0.59 0.81 ;
      RECT 0.085 0.81 0.255 2.29 ;
      RECT 4.54 2.33 8.18 2.425 ;
      RECT 5.64 2.425 8.18 2.5 ;
      RECT 7.62 1.65 7.79 2.33 ;
      RECT 8.01 2.5 8.18 2.73 ;
      RECT 7.62 1.48 8.235 1.65 ;
      RECT 8.01 2.73 8.815 2.98 ;
      RECT 7.985 0.595 8.235 1.48 ;
      RECT 4.54 2.255 6.16 2.33 ;
      RECT 5.64 2.5 5.99 2.935 ;
      RECT 5.99 1.245 6.16 2.255 ;
      RECT 5.465 1.075 6.16 1.245 ;
      RECT 5.465 0.605 5.795 1.075 ;
      RECT 3.565 2.905 4.71 3.075 ;
      RECT 4.54 2.425 4.71 2.905 ;
      RECT 3.565 2.295 3.845 2.905 ;
      RECT 3.565 0.995 3.735 2.295 ;
      RECT 3.39 0.535 3.735 0.995 ;
      RECT 8.405 2.16 8.665 2.335 ;
      RECT 7.96 1.99 8.665 2.16 ;
      RECT 7.96 1.82 8.575 1.99 ;
      RECT 8.405 0.425 8.575 1.82 ;
      RECT 7.515 0.255 9.255 0.425 ;
      RECT 7.515 0.425 7.765 1.13 ;
      RECT 9.085 0.425 9.255 0.85 ;
      RECT 9.085 0.85 10.34 1.02 ;
      RECT 9.085 1.02 9.34 1.345 ;
      RECT 10.17 0.425 10.34 0.85 ;
      RECT 10.17 0.255 11.02 0.425 ;
      RECT 10.85 0.425 11.02 0.855 ;
      RECT 10.85 0.855 11.73 1.025 ;
      RECT 11.56 1.025 11.73 1.11 ;
      RECT 11.56 1.11 13.005 1.28 ;
      RECT 11.56 1.28 11.86 1.8 ;
      RECT 12.675 1.28 13.005 1.555 ;
      RECT 13.955 2.38 14.285 2.98 ;
      RECT 13.065 2.075 14.285 2.38 ;
      RECT 14.045 1.55 14.285 2.075 ;
      RECT 14.115 0.81 14.285 1.55 ;
      RECT 13.925 0.35 14.285 0.81 ;
      RECT 0 -0.085 15.36 0.085 ;
      RECT 14.995 0.085 15.245 1.13 ;
      RECT 1.08 0.085 1.41 0.81 ;
      RECT 2.07 0.085 2.4 0.995 ;
      RECT 4.755 0.085 5.005 1.01 ;
      RECT 6.02 0.085 6.28 0.905 ;
      RECT 7.005 0.085 7.335 0.67 ;
      RECT 9.75 0.085 10 0.68 ;
      RECT 11.19 0.085 11.44 0.685 ;
      RECT 12.8 0.085 13.755 0.6 ;
      RECT 0 3.245 15.36 3.415 ;
      RECT 15.005 1.82 15.255 3.245 ;
      RECT 9.865 2.73 10.195 3.245 ;
      RECT 10.905 2.73 11.235 3.245 ;
      RECT 6.16 2.67 6.49 3.245 ;
      RECT 7.51 2.67 7.84 3.245 ;
      RECT 13.33 2.65 13.785 3.245 ;
      RECT 0.945 2.63 1.195 3.245 ;
      RECT 2.385 2.63 2.635 3.245 ;
      RECT 4.88 2.595 5.13 3.245 ;
  END
END scs8ls_sedfxtp_1

MACRO scs8ls_sedfxtp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 16.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.46 1.55 16.195 2.15 ;
        RECT 15.46 2.15 15.705 2.98 ;
        RECT 15.46 1.13 15.705 1.55 ;
        RECT 15.375 0.35 15.705 1.13 ;
    END
    ANTENNADIFFAREA 0.56 ;
  END Q

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.955 1.18 5.41 1.745 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515 1.32 1.845 1.78 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END DE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.98 0.805 1.99 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.395 1.18 6.725 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.465 1.18 4.785 1.51 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 16.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 16.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 1.58 2.725 1.75 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 1.58 15.205 1.75 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
    LAYER met1 ;
      RECT 2.495 1.735 2.785 1.78 ;
      RECT 2.495 1.595 15.265 1.735 ;
      RECT 14.975 1.735 15.265 1.78 ;
      RECT 2.495 1.55 2.785 1.595 ;
      RECT 14.975 1.55 15.265 1.595 ;
    LAYER li1 ;
      RECT 1.81 2.12 1.98 2.735 ;
      RECT 0.975 1.95 2.385 2.12 ;
      RECT 2.055 1.52 2.385 1.95 ;
      RECT 0.975 0.98 1.865 1.15 ;
      RECT 1.615 0.545 1.865 0.98 ;
      RECT 0.975 1.15 1.305 1.95 ;
      RECT 0 3.245 16.32 3.415 ;
      RECT 15.875 2.32 16.205 3.245 ;
      RECT 10.215 2.73 10.545 3.245 ;
      RECT 11.31 2.73 11.65 3.245 ;
      RECT 6.36 2.71 6.695 3.245 ;
      RECT 7.755 2.71 8.085 3.245 ;
      RECT 13.69 2.65 14.23 3.245 ;
      RECT 1.05 2.63 1.3 3.245 ;
      RECT 2.49 2.63 2.74 3.245 ;
      RECT 5.01 2.595 5.26 3.245 ;
      RECT 14.96 1.95 15.29 3.245 ;
      RECT 14.4 2.47 14.75 2.98 ;
      RECT 13.51 2.3 14.75 2.47 ;
      RECT 13.51 2.095 13.84 2.3 ;
      RECT 14.58 1.78 14.75 2.3 ;
      RECT 14.58 1.55 15.235 1.78 ;
      RECT 14.58 1.29 14.75 1.55 ;
      RECT 14.315 1.12 14.75 1.29 ;
      RECT 14.315 0.35 14.645 1.12 ;
      RECT 12.9 1.925 13.25 2.98 ;
      RECT 13.08 1.755 14.41 1.925 ;
      RECT 14.08 1.925 14.41 2.13 ;
      RECT 14.08 1.46 14.41 1.755 ;
      RECT 13.62 1.02 13.79 1.755 ;
      RECT 12.39 0.85 13.79 1.02 ;
      RECT 12.39 0.35 12.72 0.85 ;
      RECT 0 -0.085 16.32 0.085 ;
      RECT 15.875 0.085 16.205 1.13 ;
      RECT 1.055 0.085 1.385 0.81 ;
      RECT 2.045 0.085 2.375 1.005 ;
      RECT 4.885 0.085 5.215 1.01 ;
      RECT 6.235 0.085 6.495 0.68 ;
      RECT 7.235 0.085 7.485 1.13 ;
      RECT 10.1 0.085 10.365 0.68 ;
      RECT 11.635 0.085 11.885 0.68 ;
      RECT 13.21 0.085 14.145 0.68 ;
      RECT 14.875 0.085 15.205 0.95 ;
      RECT 8.645 2.2 9.005 2.35 ;
      RECT 8.205 2.02 9.005 2.2 ;
      RECT 8.205 1.82 8.815 2.02 ;
      RECT 8.645 0.425 8.815 1.82 ;
      RECT 7.665 0.255 9.495 0.425 ;
      RECT 7.665 0.425 7.995 1.13 ;
      RECT 9.325 0.425 9.495 0.85 ;
      RECT 9.325 0.85 10.705 1.02 ;
      RECT 9.325 1.02 9.655 1.345 ;
      RECT 10.535 0.425 10.705 0.85 ;
      RECT 10.535 0.255 11.465 0.425 ;
      RECT 11.295 0.425 11.465 0.85 ;
      RECT 11.295 0.85 12.21 1.02 ;
      RECT 12.04 1.02 12.21 1.19 ;
      RECT 12.04 1.19 13.45 1.36 ;
      RECT 12.04 1.36 12.37 1.8 ;
      RECT 13.12 1.36 13.45 1.585 ;
      RECT 9.715 2.39 12.73 2.56 ;
      RECT 9.715 2.35 9.885 2.39 ;
      RECT 12.56 1.755 12.73 2.39 ;
      RECT 9.525 2.02 9.885 2.35 ;
      RECT 12.56 1.53 12.91 1.755 ;
      RECT 10.75 2.05 11.125 2.22 ;
      RECT 10.955 1.52 11.125 2.05 ;
      RECT 10.955 1.36 11.8 1.52 ;
      RECT 9.915 1.19 11.8 1.36 ;
      RECT 9.915 1.36 10.245 1.49 ;
      RECT 10.875 0.595 11.125 1.19 ;
      RECT 9.185 2.52 9.545 2.98 ;
      RECT 9.185 1.83 9.355 2.52 ;
      RECT 8.985 1.66 10.785 1.83 ;
      RECT 10.455 1.53 10.785 1.66 ;
      RECT 8.985 0.595 9.155 1.66 ;
      RECT 4.67 2.37 8.425 2.425 ;
      RECT 5.8 2.425 8.425 2.52 ;
      RECT 7.865 1.65 8.035 2.37 ;
      RECT 5.8 2.52 9.015 2.54 ;
      RECT 7.865 1.48 8.475 1.65 ;
      RECT 8.255 2.54 9.015 2.69 ;
      RECT 8.225 0.595 8.475 1.48 ;
      RECT 8.765 2.69 9.015 2.98 ;
      RECT 4.67 2.255 6.225 2.37 ;
      RECT 6.055 1.065 6.225 2.255 ;
      RECT 5.8 2.54 6.13 2.935 ;
      RECT 5.675 0.895 6.225 1.065 ;
      RECT 5.675 0.605 6.005 0.895 ;
      RECT 3.67 2.905 4.84 3.075 ;
      RECT 4.67 2.425 4.84 2.905 ;
      RECT 3.67 2.295 3.95 2.905 ;
      RECT 3.67 1.005 3.84 2.295 ;
      RECT 3.51 0.545 3.84 1.005 ;
      RECT 6.895 1.53 7.615 2.2 ;
      RECT 6.895 1.01 7.065 1.53 ;
      RECT 6.675 0.35 7.065 1.01 ;
      RECT 4.01 1.915 5.885 2.085 ;
      RECT 5.62 1.415 5.885 1.915 ;
      RECT 4.125 2.255 4.5 2.735 ;
      RECT 4.01 0.605 4.715 1.01 ;
      RECT 4.125 2.085 4.295 2.255 ;
      RECT 4.01 1.01 4.295 1.915 ;
      RECT 4.01 0.255 4.295 0.605 ;
      RECT 0.085 2.29 1.64 2.46 ;
      RECT 1.47 2.46 1.64 2.905 ;
      RECT 1.47 2.905 2.32 3.075 ;
      RECT 2.15 2.46 2.32 2.905 ;
      RECT 2.15 2.29 3.5 2.46 ;
      RECT 3.25 2.46 3.5 2.975 ;
      RECT 3.33 1.345 3.5 2.29 ;
      RECT 3.17 1.175 3.5 1.345 ;
      RECT 3.17 1.005 3.34 1.175 ;
      RECT 2.865 0.675 3.34 1.005 ;
      RECT 0.085 2.46 0.51 2.98 ;
      RECT 0.085 0.35 0.565 0.81 ;
      RECT 0.085 0.81 0.255 2.29 ;
      RECT 2.555 1.515 3.07 1.845 ;
  END
END scs8ls_sedfxtp_2

MACRO scs8ls_sedfxtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 16.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.075 1.09 16.675 1.34 ;
        RECT 15.165 1.34 16.675 1.82 ;
        RECT 15.995 0.575 16.2 1.09 ;
        RECT 15.075 0.56 15.325 1.09 ;
        RECT 15.065 1.82 16.675 2.15 ;
        RECT 15.065 2.15 15.285 2.98 ;
        RECT 15.97 2.15 16.185 2.98 ;
    END
    ANTENNADIFFAREA 1.0975 ;
  END Q

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.955 1.18 5.37 1.745 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535 1.32 1.865 1.78 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END DE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.98 0.825 1.99 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.455 1.18 7.075 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.18 4.785 1.51 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 16.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 16.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 1.58 2.725 1.75 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 1.58 14.725 1.75 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
    LAYER met1 ;
      RECT 2.495 1.735 2.785 1.78 ;
      RECT 2.495 1.595 14.785 1.735 ;
      RECT 14.495 1.735 14.785 1.78 ;
      RECT 2.495 1.55 2.785 1.595 ;
      RECT 14.495 1.55 14.785 1.595 ;
    LAYER li1 ;
      RECT 3.995 1.915 5.86 2.085 ;
      RECT 5.58 1.415 5.86 1.915 ;
      RECT 4.105 2.255 4.46 2.735 ;
      RECT 3.995 0.605 4.585 1.01 ;
      RECT 4.105 2.085 4.275 2.255 ;
      RECT 3.995 1.01 4.275 1.915 ;
      RECT 3.995 0.255 4.275 0.605 ;
      RECT 0.085 2.29 1.625 2.46 ;
      RECT 1.455 2.46 1.625 2.905 ;
      RECT 1.455 2.905 2.305 3.075 ;
      RECT 2.135 2.46 2.305 2.905 ;
      RECT 2.135 2.29 3.485 2.46 ;
      RECT 3.235 2.46 3.485 2.975 ;
      RECT 3.315 1.345 3.485 2.29 ;
      RECT 2.85 1.175 3.485 1.345 ;
      RECT 2.85 0.545 3.18 1.175 ;
      RECT 0.085 2.46 0.495 2.98 ;
      RECT 0.085 0.34 0.55 0.81 ;
      RECT 0.085 0.81 0.255 2.29 ;
      RECT 2.535 1.52 3.055 1.85 ;
      RECT 1.795 2.12 1.965 2.735 ;
      RECT 0.995 1.95 2.365 2.12 ;
      RECT 2.115 1.52 2.365 1.95 ;
      RECT 0.995 0.98 1.85 1.15 ;
      RECT 1.6 0.545 1.85 0.98 ;
      RECT 0.995 1.15 1.325 1.95 ;
      RECT 0 3.245 16.8 3.415 ;
      RECT 16.365 2.32 16.695 3.245 ;
      RECT 9.96 2.73 10.29 3.245 ;
      RECT 10.995 2.73 11.325 3.245 ;
      RECT 6.26 2.675 6.59 3.245 ;
      RECT 7.61 2.675 7.94 3.245 ;
      RECT 13.335 2.65 13.875 3.245 ;
      RECT 1.035 2.63 1.285 3.245 ;
      RECT 2.475 2.63 2.725 3.245 ;
      RECT 4.97 2.595 5.22 3.245 ;
      RECT 14.565 1.95 14.895 3.245 ;
      RECT 15.465 2.32 15.795 3.245 ;
      RECT 0 -0.085 16.8 0.085 ;
      RECT 16.37 0.085 16.7 0.92 ;
      RECT 7.095 0.085 7.425 0.67 ;
      RECT 9.84 0.085 10.09 0.69 ;
      RECT 11.28 0.085 11.53 0.69 ;
      RECT 12.855 0.085 13.835 0.68 ;
      RECT 14.565 0.085 14.895 1.34 ;
      RECT 15.495 0.085 15.825 0.92 ;
      RECT 4.765 0.085 5.095 1.01 ;
      RECT 6.11 0.085 6.36 0.905 ;
      RECT 2.03 0.085 2.36 1.005 ;
      RECT 1.04 0.085 1.37 0.81 ;
      RECT 14.045 2.35 14.395 2.98 ;
      RECT 13.155 2.18 14.395 2.35 ;
      RECT 13.155 2.095 13.485 2.18 ;
      RECT 14.225 1.78 14.395 2.18 ;
      RECT 14.225 1.55 14.755 1.78 ;
      RECT 14.225 0.81 14.395 1.55 ;
      RECT 14.005 0.35 14.395 0.81 ;
      RECT 12.465 1.925 12.895 2.98 ;
      RECT 12.725 1.755 14.055 1.925 ;
      RECT 13.725 1.925 14.055 1.99 ;
      RECT 13.265 1.02 14.055 1.755 ;
      RECT 12.035 0.99 14.055 1.02 ;
      RECT 13.725 0.98 14.055 0.99 ;
      RECT 12.035 0.85 13.435 0.99 ;
      RECT 12.035 0.35 12.365 0.85 ;
      RECT 8.495 2.165 8.83 2.335 ;
      RECT 8.06 1.995 8.83 2.165 ;
      RECT 8.06 1.82 8.665 1.995 ;
      RECT 8.495 0.425 8.665 1.82 ;
      RECT 7.605 0.255 9.505 0.425 ;
      RECT 7.605 0.425 7.855 1.13 ;
      RECT 9.175 0.425 9.505 0.86 ;
      RECT 9.175 0.86 10.43 1.03 ;
      RECT 9.175 1.03 9.505 1.255 ;
      RECT 10.26 0.425 10.43 0.86 ;
      RECT 10.26 0.255 11.11 0.425 ;
      RECT 10.94 0.425 11.11 0.86 ;
      RECT 10.94 0.86 11.855 1.03 ;
      RECT 11.685 1.03 11.855 1.19 ;
      RECT 11.685 1.19 13.095 1.36 ;
      RECT 11.685 1.36 11.955 1.8 ;
      RECT 12.765 1.36 13.095 1.585 ;
      RECT 9.53 2.39 12.295 2.56 ;
      RECT 9.53 2.33 9.7 2.39 ;
      RECT 12.125 1.755 12.295 2.39 ;
      RECT 9.34 2 9.7 2.33 ;
      RECT 12.125 1.53 12.555 1.755 ;
      RECT 10.475 1.97 10.925 2.22 ;
      RECT 10.755 1.53 10.925 1.97 ;
      RECT 10.755 1.37 11.475 1.53 ;
      RECT 9.715 1.2 11.475 1.37 ;
      RECT 9.715 1.37 10.045 1.405 ;
      RECT 10.6 0.595 10.77 1.2 ;
      RECT 9 2.52 9.36 2.98 ;
      RECT 9 1.8 9.17 2.52 ;
      RECT 8.835 1.63 10.585 1.8 ;
      RECT 10.255 1.54 10.585 1.63 ;
      RECT 8.835 0.595 9.005 1.63 ;
      RECT 4.63 2.335 8.325 2.425 ;
      RECT 5.73 2.425 8.325 2.505 ;
      RECT 7.72 1.65 7.89 2.335 ;
      RECT 8.155 2.505 8.83 2.98 ;
      RECT 7.72 1.48 8.325 1.65 ;
      RECT 8.075 0.595 8.325 1.48 ;
      RECT 4.63 2.255 6.2 2.335 ;
      RECT 5.73 2.505 6.06 2.935 ;
      RECT 6.03 1.245 6.2 2.255 ;
      RECT 5.555 1.075 6.2 1.245 ;
      RECT 5.555 0.605 5.885 1.075 ;
      RECT 3.655 2.905 4.8 3.075 ;
      RECT 4.63 2.425 4.8 2.905 ;
      RECT 3.655 2.295 3.935 2.905 ;
      RECT 3.655 1.005 3.825 2.295 ;
      RECT 3.35 0.675 3.825 1.005 ;
      RECT 6.71 1.785 7.49 2.165 ;
      RECT 7.245 1.01 7.415 1.785 ;
      RECT 6.54 0.84 7.415 1.01 ;
      RECT 6.54 0.35 6.87 0.84 ;
  END
END scs8ls_sedfxtp_4

MACRO scs8ls_tap_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.48 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.89 0.39 3.065 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.265 0.39 1.44 ;
    END
  END vnb

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.48 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.48 3.575 ;
    END
  END vpwr
  OBS
    LAYER li1 ;
      RECT 0 -0.085 0.48 0.085 ;
      RECT 0 3.245 0.48 3.415 ;
    LAYER mcon ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_tap_1

MACRO scs8ls_tap_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.89 0.87 3.065 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.265 0.87 1.44 ;
    END
  END vnb

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.96 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.96 3.575 ;
    END
  END vpwr
  OBS
    LAYER li1 ;
      RECT 0 -0.085 0.96 0.085 ;
      RECT 0 3.245 0.96 3.415 ;
    LAYER mcon ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_tap_2

MACRO scs8ls_tapvgnd2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.48 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.48 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.48 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.08 2.275 0.4 2.535 ;
    END
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb
  OBS
    LAYER li1 ;
      RECT 0 3.245 0.48 3.415 ;
      RECT 0.09 0.085 0.39 1.44 ;
      RECT 0 -0.085 0.48 0.085 ;
      RECT 0.09 1.89 0.39 3.065 ;
    LAYER mcon ;
      RECT 0.155 2.32 0.325 2.49 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_tapvgnd2_1

MACRO scs8ls_tapvgnd_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.48 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.48 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.48 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.08 2.645 0.4 2.905 ;
    END
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb
  OBS
    LAYER li1 ;
      RECT 0 3.245 0.48 3.415 ;
      RECT 0.09 0.085 0.39 1.44 ;
      RECT 0 -0.085 0.48 0.085 ;
      RECT 0.09 1.89 0.39 3.065 ;
    LAYER mcon ;
      RECT 0.155 2.69 0.325 2.86 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_tapvgnd_1

MACRO scs8ls_tapvpwrvgnd_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.48 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.48 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.48 3.575 ;
    END
  END vpwr
  OBS
    LAYER li1 ;
      RECT 0 3.245 0.48 3.415 ;
      RECT 0.09 2.205 0.39 3.245 ;
      RECT 0.09 0.085 0.39 1.105 ;
      RECT 0 -0.085 0.48 0.085 ;
    LAYER mcon ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_tapvpwrvgnd_1

MACRO scs8ls_xnor2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 1.435 1.345 1.78 ;
        RECT 1.175 1.78 1.345 1.95 ;
        RECT 1.175 1.95 2.185 2.12 ;
        RECT 2.015 1.68 2.185 1.95 ;
        RECT 2.015 1.35 2.465 1.68 ;
    END
    ANTENNAGATEAREA 0.501 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 2.29 2.685 2.98 ;
        RECT 2.355 2.02 2.685 2.29 ;
        RECT 2.355 1.85 3.275 2.02 ;
        RECT 3.105 1.13 3.275 1.85 ;
        RECT 2.975 0.35 3.275 1.13 ;
    END
    ANTENNADIFFAREA 0.6998 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515 1.35 1.845 1.78 ;
    END
    ANTENNAGATEAREA 0.501 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.855 2.19 3.185 3.245 ;
      RECT 0.175 2.29 0.505 3.245 ;
      RECT 0.175 1.905 0.425 2.29 ;
      RECT 1.415 2.29 1.745 3.245 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 0.105 0.085 0.435 1.255 ;
      RECT 1.935 0.085 2.265 0.5 ;
      RECT 0.605 1.085 2.805 1.18 ;
      RECT 2.635 1.18 2.805 1.3 ;
      RECT 0.895 1.01 2.805 1.085 ;
      RECT 2.635 1.3 2.935 1.63 ;
      RECT 0.605 1.255 0.775 1.95 ;
      RECT 0.675 2.12 1.005 2.785 ;
      RECT 0.605 1.95 1.005 2.12 ;
      RECT 0.605 1.18 1.225 1.255 ;
      RECT 0.895 0.575 1.225 1.01 ;
      RECT 1.435 0.67 2.77 0.84 ;
      RECT 1.435 0.51 1.765 0.67 ;
      RECT 2.44 0.51 2.77 0.67 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_xnor2_1

MACRO scs8ls_xnor2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.35 4.855 1.68 ;
        RECT 4.445 1.68 4.675 1.72 ;
        RECT 3.025 1.72 4.675 1.89 ;
        RECT 3.025 1.55 3.355 1.72 ;
        RECT 3.005 1.18 3.355 1.55 ;
    END
    ANTENNAGATEAREA 0.819 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.107 LAYER met1 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.925 1.18 4.255 1.55 ;
        RECT 3.925 1.01 5.195 1.18 ;
        RECT 5.025 1.18 5.195 2.06 ;
        RECT 2.605 2.06 5.195 2.23 ;
        RECT 2.605 1.89 2.775 2.06 ;
        RECT 1.345 1.72 2.775 1.89 ;
        RECT 1.345 1.35 1.675 1.72 ;
    END
    ANTENNAGATEAREA 0.819 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 2.4 4.135 2.49 ;
        RECT 2.045 2.49 4.135 2.57 ;
        RECT 0.085 2.32 2.435 2.4 ;
        RECT 2.045 2.06 2.435 2.32 ;
        RECT 2.045 2.57 2.435 2.98 ;
        RECT 3.805 2.57 4.135 2.735 ;
        RECT 0.085 1.01 0.255 2.32 ;
        RECT 0.085 0.84 0.835 1.01 ;
        RECT 0.665 0.425 0.835 0.84 ;
        RECT 0.665 0.255 2.575 0.425 ;
        RECT 2.19 0.425 2.575 0.5 ;
    END
    ANTENNADIFFAREA 1.0728 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 0.575 1.365 0.865 1.41 ;
      RECT 0.575 1.225 3.265 1.365 ;
      RECT 2.975 1.365 3.265 1.41 ;
      RECT 0.575 1.18 0.865 1.225 ;
      RECT 2.975 1.18 3.265 1.225 ;
    LAYER li1 ;
      RECT 0 -0.085 5.28 0.085 ;
      RECT 3.265 0.085 3.6 0.5 ;
      RECT 4.31 0.085 4.655 0.5 ;
      RECT 0.115 0.085 0.495 0.67 ;
      RECT 0 3.245 5.28 3.415 ;
      RECT 4.805 2.4 5.135 3.245 ;
      RECT 0.115 2.66 0.445 3.245 ;
      RECT 1.23 2.66 1.875 3.245 ;
      RECT 2.64 2.74 2.97 3.245 ;
      RECT 3.26 2.905 4.635 3.075 ;
      RECT 4.305 2.4 4.635 2.905 ;
      RECT 3.26 2.74 3.6 2.905 ;
      RECT 2.755 0.84 3.085 1.01 ;
      RECT 1.68 0.67 5.165 0.84 ;
      RECT 3.78 0.49 4.11 0.67 ;
      RECT 4.835 0.49 5.165 0.67 ;
      RECT 2.755 0.35 3.085 0.67 ;
      RECT 1.68 0.595 2.01 0.67 ;
      RECT 1.005 1.01 2.585 1.18 ;
      RECT 1.915 1.18 2.585 1.55 ;
      RECT 1.005 0.635 1.45 1.01 ;
      RECT 0.65 1.82 1.175 2.15 ;
      RECT 1.005 1.18 1.175 1.82 ;
      RECT 0.425 1.18 0.835 1.55 ;
    LAYER mcon ;
      RECT 3.035 1.21 3.205 1.38 ;
      RECT 0.635 1.21 0.805 1.38 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_xnor2_2

MACRO scs8ls_xnor2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.35 5.835 1.775 ;
    END
    ANTENNAGATEAREA 1.56 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.779 LAYER met1 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.35 8.155 1.765 ;
        RECT 6.365 1.765 6.535 1.945 ;
        RECT 1.985 1.945 6.535 2.115 ;
        RECT 1.985 1.68 2.155 1.945 ;
        RECT 1.485 1.35 2.155 1.68 ;
    END
    ANTENNAGATEAREA 1.56 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.325 1.935 8.555 2.105 ;
        RECT 7.325 2.105 7.655 2.285 ;
        RECT 8.225 2.105 8.555 2.735 ;
        RECT 8.325 1.18 8.495 1.935 ;
        RECT 2.545 2.285 7.655 2.455 ;
        RECT 3.035 1.01 8.495 1.18 ;
        RECT 7.325 2.455 7.655 2.735 ;
        RECT 3.035 0.595 3.365 1.01 ;
        RECT 4.06 0.595 4.39 1.01 ;
    END
    ANTENNADIFFAREA 1.4742 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 1.055 1.735 1.345 1.78 ;
      RECT 1.055 1.595 4.705 1.735 ;
      RECT 4.415 1.735 4.705 1.78 ;
      RECT 1.055 1.55 1.345 1.595 ;
      RECT 4.415 1.55 4.705 1.595 ;
    LAYER li1 ;
      RECT 0.115 0.98 1.375 1.15 ;
      RECT 1.045 0.6 1.375 0.98 ;
      RECT 0.115 0.35 0.365 0.98 ;
      RECT 1.045 0.35 2.305 0.6 ;
      RECT 1.085 1.65 1.315 1.78 ;
      RECT 0.545 1.32 1.315 1.65 ;
      RECT 2.395 1.35 4.085 1.68 ;
      RECT 2.395 1.18 2.565 1.35 ;
      RECT 1.545 1.01 2.565 1.18 ;
      RECT 1.545 0.77 1.875 1.01 ;
      RECT 8.675 0.84 9.005 1.13 ;
      RECT 4.56 0.67 9.005 0.84 ;
      RECT 4.56 0.425 4.89 0.67 ;
      RECT 5.58 0.35 5.91 0.67 ;
      RECT 6.6 0.35 6.93 0.67 ;
      RECT 7.655 0.35 7.985 0.67 ;
      RECT 8.675 0.35 9.005 0.67 ;
      RECT 2.535 0.255 4.89 0.425 ;
      RECT 2.535 0.425 2.865 0.84 ;
      RECT 3.535 0.425 3.865 0.84 ;
      RECT 3.58 2.795 4.59 2.955 ;
      RECT 1.465 2.625 4.59 2.795 ;
      RECT 1.465 2.12 1.795 2.625 ;
      RECT 0.565 1.95 1.795 2.12 ;
      RECT 0.565 2.12 0.895 2.7 ;
      RECT 0.565 1.82 0.895 1.95 ;
      RECT 6.875 2.905 9.005 3.075 ;
      RECT 8.755 1.935 9.005 2.905 ;
      RECT 4.81 2.625 7.125 2.795 ;
      RECT 6.875 2.795 7.125 2.905 ;
      RECT 4.81 2.795 5.06 2.98 ;
      RECT 5.805 2.795 6.135 2.98 ;
      RECT 7.855 2.275 8.025 2.905 ;
      RECT 0 3.245 9.12 3.415 ;
      RECT 1.095 2.29 1.265 3.245 ;
      RECT 0.115 1.82 0.365 3.245 ;
      RECT 2 2.965 2.34 3.245 ;
      RECT 6.34 2.965 6.67 3.245 ;
      RECT 3.08 2.965 3.41 3.245 ;
      RECT 5.265 2.965 5.6 3.245 ;
      RECT 0 -0.085 9.12 0.085 ;
      RECT 5.07 0.085 5.4 0.5 ;
      RECT 6.09 0.085 6.42 0.5 ;
      RECT 7.11 0.085 7.475 0.5 ;
      RECT 8.165 0.085 8.495 0.5 ;
      RECT 0.545 0.085 0.875 0.81 ;
    LAYER mcon ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 1.115 1.58 1.285 1.75 ;
      RECT 4.475 1.58 4.645 1.75 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
  END
END scs8ls_xnor2_4

MACRO scs8ls_xnor3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845 1.425 7.205 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995 1.35 1.325 1.78 ;
    END
    ANTENNAGATEAREA 0.381 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.705 1.35 4.375 1.78 ;
    END
    ANTENNAGATEAREA 0.693 ;
  END B

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.44 0.445 1.17 ;
        RECT 0.085 1.17 0.255 1.84 ;
        RECT 0.085 1.84 0.355 2.98 ;
    END
    ANTENNADIFFAREA 0.5301 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 2.015 1.365 2.305 1.41 ;
      RECT 2.015 1.225 5.665 1.365 ;
      RECT 5.375 1.365 5.665 1.41 ;
      RECT 2.015 1.18 2.305 1.225 ;
      RECT 5.375 1.18 5.665 1.225 ;
      RECT 5.855 1.365 6.145 1.41 ;
      RECT 5.855 1.225 8.065 1.365 ;
      RECT 7.775 1.365 8.065 1.41 ;
      RECT 5.855 1.18 6.145 1.225 ;
      RECT 7.775 1.18 8.065 1.225 ;
    LAYER li1 ;
      RECT 3.92 1.95 4.715 2.2 ;
      RECT 4.545 1.685 4.715 1.95 ;
      RECT 4.545 1.355 5.045 1.685 ;
      RECT 4.545 1.18 4.715 1.355 ;
      RECT 3.905 1.01 4.715 1.18 ;
      RECT 1.315 1.95 1.665 2.5 ;
      RECT 1.495 1.75 1.665 1.95 ;
      RECT 1.495 1.58 2.845 1.75 ;
      RECT 2.515 1.75 2.845 1.81 ;
      RECT 2.515 1.48 2.845 1.58 ;
      RECT 1.495 1.17 1.665 1.58 ;
      RECT 1.135 1 1.665 1.17 ;
      RECT 2.85 2.03 3.185 2.2 ;
      RECT 3.015 1.31 3.185 2.03 ;
      RECT 1.835 1.14 3.185 1.31 ;
      RECT 1.835 1.31 2.275 1.41 ;
      RECT 1.835 0.595 2.165 1.14 ;
      RECT 0.975 2.905 2.655 3.075 ;
      RECT 2.325 2.71 2.655 2.905 ;
      RECT 0.975 2.12 1.145 2.905 ;
      RECT 0.615 1.95 1.145 2.12 ;
      RECT 0.615 0.66 1.665 0.83 ;
      RECT 1.495 0.425 1.665 0.66 ;
      RECT 1.495 0.255 2.665 0.425 ;
      RECT 2.335 0.425 2.665 0.97 ;
      RECT 0.615 1.67 0.785 1.95 ;
      RECT 0.425 1.34 0.785 1.67 ;
      RECT 0.615 0.83 0.785 1.34 ;
      RECT 6.08 1.935 6.25 2.395 ;
      RECT 5.435 1.765 6.25 1.935 ;
      RECT 5.435 1.41 5.605 1.765 ;
      RECT 5.315 1.185 5.605 1.41 ;
      RECT 5.02 1.18 5.605 1.185 ;
      RECT 5.02 1.015 5.485 1.18 ;
      RECT 5.55 2.565 6.59 2.735 ;
      RECT 5.55 2.105 5.88 2.565 ;
      RECT 6.42 1.595 6.59 2.565 ;
      RECT 5.775 1.425 6.59 1.595 ;
      RECT 5.775 0.935 6.085 1.425 ;
      RECT 7.79 2.19 8.075 2.93 ;
      RECT 7.835 1.255 8.075 2.19 ;
      RECT 7.795 0.585 8.075 1.255 ;
      RECT 4.49 2.905 7.09 3.075 ;
      RECT 6.76 2.12 7.09 2.905 ;
      RECT 6.76 1.95 7.62 2.12 ;
      RECT 7.415 1.755 7.62 1.95 ;
      RECT 7.415 1.425 7.665 1.755 ;
      RECT 7.415 1.255 7.62 1.425 ;
      RECT 6.705 1.085 7.62 1.255 ;
      RECT 6.705 0.425 7.035 1.085 ;
      RECT 4.465 0.255 7.035 0.425 ;
      RECT 4.49 2.71 4.82 2.905 ;
      RECT 4.465 0.425 4.84 0.5 ;
      RECT 1.875 2.37 5.265 2.54 ;
      RECT 5.015 2.54 5.265 2.575 ;
      RECT 5.015 1.855 5.265 2.37 ;
      RECT 2.835 0.765 5.18 0.84 ;
      RECT 2.835 0.67 6.535 0.765 ;
      RECT 6.255 0.765 6.535 1.21 ;
      RECT 5.01 0.595 6.535 0.67 ;
      RECT 1.875 2.54 2.125 2.735 ;
      RECT 1.875 1.95 2.125 2.37 ;
      RECT 3.355 0.97 3.525 2.37 ;
      RECT 2.835 0.84 3.525 0.97 ;
      RECT 2.835 0.35 3.165 0.67 ;
      RECT 0.625 0.085 0.955 0.49 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 3.395 0.085 3.725 0.5 ;
      RECT 7.205 0.085 7.615 0.915 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 3.395 2.71 3.725 3.245 ;
      RECT 0.555 2.29 0.805 3.245 ;
      RECT 7.26 2.29 7.59 3.245 ;
    LAYER mcon ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 1.21 5.605 1.38 ;
      RECT 5.915 1.21 6.085 1.38 ;
      RECT 2.075 1.21 2.245 1.38 ;
      RECT 7.835 1.21 8.005 1.38 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
  END
END scs8ls_xnor3_1

MACRO scs8ls_xnor3_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955 1.375 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845 1.35 7.175 1.78 ;
    END
    ANTENNAGATEAREA 0.381 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.735 1.35 4.405 1.78 ;
    END
    ANTENNAGATEAREA 0.693 ;
  END B

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.765 0.44 8.095 1.17 ;
        RECT 7.925 1.17 8.095 1.84 ;
        RECT 7.75 1.84 8.095 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 2.495 1.365 2.785 1.41 ;
      RECT 2.495 1.225 5.185 1.365 ;
      RECT 4.895 1.365 5.185 1.41 ;
      RECT 2.495 1.18 2.785 1.225 ;
      RECT 4.895 1.18 5.185 1.225 ;
      RECT 0.095 1.365 0.385 1.41 ;
      RECT 0.095 1.225 1.825 1.365 ;
      RECT 1.535 1.365 1.825 1.41 ;
      RECT 0.095 1.18 0.385 1.225 ;
      RECT 1.535 1.18 1.825 1.225 ;
    LAYER li1 ;
      RECT 6.07 2.565 6.32 2.735 ;
      RECT 4.585 2.54 6.32 2.565 ;
      RECT 2.835 2.395 6.32 2.54 ;
      RECT 2.835 2.37 4.755 2.395 ;
      RECT 6.07 1.975 6.32 2.395 ;
      RECT 4.585 0.965 4.755 2.37 ;
      RECT 4.585 0.785 5.16 0.965 ;
      RECT 2.555 0.765 5.16 0.785 ;
      RECT 1.625 0.615 5.16 0.765 ;
      RECT 4.83 0.35 5.16 0.615 ;
      RECT 2.835 2.54 3.065 2.62 ;
      RECT 2.835 1.875 3.145 2.37 ;
      RECT 1.625 0.765 1.955 0.995 ;
      RECT 1.625 0.595 2.725 0.615 ;
      RECT 3.395 1.95 4.255 2.2 ;
      RECT 3.395 0.955 4.09 1.125 ;
      RECT 3.395 1.705 3.565 1.95 ;
      RECT 3.155 1.375 3.565 1.705 ;
      RECT 3.395 1.125 3.565 1.375 ;
      RECT 6.505 1.95 6.87 2.5 ;
      RECT 6.505 1.805 6.675 1.95 ;
      RECT 5.325 1.475 6.675 1.805 ;
      RECT 6.39 1.17 6.675 1.475 ;
      RECT 6.39 1 6.72 1.17 ;
      RECT 4.925 1.975 5.335 2.225 ;
      RECT 4.925 1.305 5.155 1.975 ;
      RECT 4.925 1.135 6.16 1.305 ;
      RECT 5.83 0.595 6.16 1.135 ;
      RECT 1.885 1.72 2.105 2.395 ;
      RECT 1.885 1.55 2.755 1.72 ;
      RECT 2.555 1.285 2.755 1.55 ;
      RECT 2.555 0.955 2.985 1.285 ;
      RECT 7.41 1.34 7.755 1.67 ;
      RECT 5.535 2.905 7.21 3.075 ;
      RECT 7.04 2.12 7.21 2.905 ;
      RECT 7.04 1.95 7.58 2.12 ;
      RECT 7.41 1.67 7.58 1.95 ;
      RECT 7.41 1.18 7.58 1.34 ;
      RECT 6.89 1.01 7.58 1.18 ;
      RECT 6.89 0.83 7.06 1.01 ;
      RECT 6.33 0.66 7.06 0.83 ;
      RECT 5.535 2.735 5.865 2.905 ;
      RECT 6.33 0.425 6.5 0.66 ;
      RECT 5.33 0.255 6.5 0.425 ;
      RECT 5.33 0.425 5.66 0.965 ;
      RECT 1.545 2.565 2.605 2.735 ;
      RECT 2.275 1.89 2.605 2.565 ;
      RECT 1.545 1.38 1.715 2.565 ;
      RECT 1.545 1.165 2.385 1.38 ;
      RECT 2.135 0.935 2.385 1.165 ;
      RECT 0.085 2.29 0.445 2.885 ;
      RECT 0.085 1.065 0.325 2.29 ;
      RECT 0.085 0.385 0.405 1.065 ;
      RECT 1.095 2.905 3.675 3.075 ;
      RECT 3.345 2.71 3.675 2.905 ;
      RECT 1.095 2.12 1.375 2.905 ;
      RECT 0.495 1.95 1.375 2.12 ;
      RECT 0.575 1.035 1.345 1.205 ;
      RECT 1.095 0.425 1.345 1.035 ;
      RECT 1.095 0.255 3.53 0.425 ;
      RECT 3.2 0.425 3.53 0.445 ;
      RECT 0.495 1.235 0.745 1.95 ;
      RECT 0.575 1.205 0.745 1.235 ;
      RECT 0 -0.085 8.64 0.085 ;
      RECT 8.275 0.085 8.525 1.25 ;
      RECT 7.23 0.49 7.585 0.84 ;
      RECT 6.9 0.085 7.585 0.49 ;
      RECT 0.585 0.085 0.915 0.865 ;
      RECT 4.27 0.085 4.6 0.445 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 8.28 1.82 8.53 3.245 ;
      RECT 4.455 2.735 4.785 3.245 ;
      RECT 0.645 2.305 0.925 3.245 ;
      RECT 7.38 2.29 7.55 3.245 ;
    LAYER mcon ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.555 1.21 2.725 1.38 ;
      RECT 1.595 1.21 1.765 1.38 ;
      RECT 4.955 1.21 5.125 1.38 ;
      RECT 0.155 1.21 0.325 1.38 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_xnor3_2

MACRO scs8ls_xnor3_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.915 1.375 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.78 1.35 7.11 1.78 ;
    END
    ANTENNAGATEAREA 0.381 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.94 1.35 4.27 1.78 ;
    END
    ANTENNAGATEAREA 0.693 ;
  END B

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.205 0.44 9.535 1.42 ;
        RECT 8.47 1.42 9.535 1.625 ;
        RECT 9.18 1.625 9.535 2.98 ;
        RECT 8.47 1.625 8.64 1.84 ;
        RECT 8.47 1.17 8.675 1.42 ;
        RECT 8.28 1.84 8.64 2.98 ;
        RECT 8.345 0.47 8.675 1.17 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 1.95 1.765 2.12 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 1.95 0.325 2.12 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 1.95 5.125 2.12 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 1.95 2.245 2.12 ;
    LAYER met1 ;
      RECT 2.015 2.105 2.305 2.15 ;
      RECT 2.015 1.965 5.185 2.105 ;
      RECT 4.895 2.105 5.185 2.15 ;
      RECT 2.015 1.92 2.305 1.965 ;
      RECT 4.895 1.92 5.185 1.965 ;
      RECT 0.095 2.105 0.385 2.15 ;
      RECT 0.095 1.965 1.825 2.105 ;
      RECT 1.535 2.105 1.825 2.15 ;
      RECT 0.095 1.92 0.385 1.965 ;
      RECT 1.535 1.92 1.825 1.965 ;
    LAYER li1 ;
      RECT 6.02 2.56 6.27 2.735 ;
      RECT 4.44 2.54 6.27 2.56 ;
      RECT 2.895 2.39 6.27 2.54 ;
      RECT 2.895 2.37 4.61 2.39 ;
      RECT 6.02 1.97 6.27 2.39 ;
      RECT 4.44 1.03 4.61 2.37 ;
      RECT 4.44 0.785 5.16 1.03 ;
      RECT 2.555 0.765 5.16 0.785 ;
      RECT 1.625 0.615 5.16 0.765 ;
      RECT 4.83 0.35 5.16 0.615 ;
      RECT 2.895 2.54 3.145 2.545 ;
      RECT 2.895 1.875 3.145 2.37 ;
      RECT 1.625 0.765 1.955 0.995 ;
      RECT 1.625 0.595 2.725 0.615 ;
      RECT 7.32 1.34 8.3 1.67 ;
      RECT 5.485 2.905 7.315 3.075 ;
      RECT 7.13 2.12 7.315 2.905 ;
      RECT 7.13 1.95 7.49 2.12 ;
      RECT 7.32 1.67 7.49 1.95 ;
      RECT 7.32 1.18 7.49 1.34 ;
      RECT 6.89 1.01 7.49 1.18 ;
      RECT 6.89 0.83 7.06 1.01 ;
      RECT 6.33 0.66 7.06 0.83 ;
      RECT 5.485 2.73 5.815 2.905 ;
      RECT 6.33 0.425 6.5 0.66 ;
      RECT 5.33 0.255 6.5 0.425 ;
      RECT 5.33 0.425 5.66 1.01 ;
      RECT 0 3.245 10.08 3.415 ;
      RECT 9.71 1.82 9.96 3.245 ;
      RECT 4.39 2.73 4.72 3.245 ;
      RECT 0.565 2.29 0.895 3.245 ;
      RECT 7.485 2.29 8.11 3.245 ;
      RECT 7.685 1.84 8.11 2.29 ;
      RECT 8.81 1.82 8.98 3.245 ;
      RECT 0 -0.085 10.08 0.085 ;
      RECT 9.715 0.085 9.965 1.25 ;
      RECT 7.915 0.84 8.165 1.17 ;
      RECT 7.23 0.49 8.165 0.84 ;
      RECT 6.9 0.085 8.165 0.49 ;
      RECT 0.665 0.085 0.995 0.865 ;
      RECT 4.27 0.085 4.6 0.445 ;
      RECT 8.855 0.085 9.025 1.25 ;
      RECT 4.78 1.95 5.28 2.22 ;
      RECT 4.78 1.38 4.95 1.95 ;
      RECT 4.78 1.21 6.16 1.38 ;
      RECT 5.405 1.18 6.16 1.21 ;
      RECT 5.83 0.595 6.16 1.18 ;
      RECT 3.6 1.95 4.27 2.2 ;
      RECT 3.6 0.955 4.09 1.125 ;
      RECT 3.6 1.705 3.77 1.95 ;
      RECT 2.995 1.375 3.77 1.705 ;
      RECT 3.6 1.125 3.77 1.375 ;
      RECT 1.065 2.905 3.68 3.075 ;
      RECT 3.35 2.71 3.68 2.905 ;
      RECT 1.065 2.12 1.395 2.905 ;
      RECT 0.535 1.95 1.395 2.12 ;
      RECT 0.455 1.035 1.425 1.205 ;
      RECT 1.175 0.425 1.425 1.035 ;
      RECT 1.175 0.255 3.53 0.425 ;
      RECT 3.2 0.425 3.53 0.445 ;
      RECT 0.535 1.465 0.705 1.95 ;
      RECT 0.455 1.205 0.705 1.465 ;
      RECT 1.935 2.12 2.135 2.155 ;
      RECT 1.935 1.675 2.245 2.12 ;
      RECT 1.935 1.505 2.755 1.675 ;
      RECT 2.555 1.205 2.755 1.505 ;
      RECT 2.555 0.955 3.02 1.205 ;
      RECT 1.565 2.565 2.725 2.735 ;
      RECT 2.305 2.29 2.725 2.565 ;
      RECT 1.565 1.375 1.765 2.565 ;
      RECT 1.595 1.335 1.765 1.375 ;
      RECT 1.595 1.165 2.385 1.335 ;
      RECT 2.135 0.935 2.385 1.165 ;
      RECT 6.44 1.99 6.96 2.5 ;
      RECT 6.44 1.72 6.61 1.99 ;
      RECT 5.12 1.55 6.61 1.72 ;
      RECT 5.12 1.72 5.45 1.78 ;
      RECT 6.39 1.17 6.61 1.55 ;
      RECT 6.39 1 6.72 1.17 ;
      RECT 0.085 1.845 0.365 2.885 ;
      RECT 0.085 0.865 0.285 1.845 ;
      RECT 0.085 0.365 0.495 0.865 ;
  END
END scs8ls_xnor3_4

MACRO scs8ls_xor2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 0.415 2.97 0.98 ;
        RECT 2.525 0.98 3.755 1.15 ;
        RECT 3.585 1.15 3.755 1.82 ;
        RECT 3.365 1.82 3.755 2.98 ;
    END
    ANTENNADIFFAREA 0.6972 ;
  END X

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.285 1.365 2.845 1.695 ;
        RECT 2.515 1.695 2.845 1.78 ;
        RECT 2.515 1.35 2.845 1.365 ;
    END
    ANTENNAGATEAREA 0.512 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.775 1.615 ;
    END
    ANTENNAGATEAREA 0.512 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.755 2.46 2.085 2.98 ;
      RECT 1.755 2.29 3.195 2.46 ;
      RECT 2.865 2.46 3.195 2.98 ;
      RECT 3.025 1.32 3.415 1.65 ;
      RECT 0.945 1.95 3.195 2.12 ;
      RECT 3.025 1.65 3.195 1.95 ;
      RECT 0.945 1.04 1.115 1.95 ;
      RECT 0.945 2.12 1.525 2.98 ;
      RECT 0.945 0.71 1.64 1.04 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 2.255 2.65 2.695 3.245 ;
      RECT 0.325 1.94 0.655 3.245 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 0.175 0.085 0.775 0.99 ;
      RECT 1.82 0.085 2.15 1.195 ;
      RECT 3.21 0.085 3.54 0.745 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_xor2_1

MACRO scs8ls_xor2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.355 0.35 4.685 0.67 ;
        RECT 3.33 0.67 4.685 0.84 ;
        RECT 4.355 0.84 4.685 1.85 ;
        RECT 3.33 0.595 3.66 0.67 ;
        RECT 3.025 1.85 4.685 2.02 ;
        RECT 3.025 2.02 3.195 2.735 ;
    END
    ANTENNADIFFAREA 0.7541 ;
  END X

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.18 4.145 1.55 ;
        RECT 1.155 1.01 4.145 1.18 ;
        RECT 1.155 1.18 1.485 1.45 ;
    END
    ANTENNAGATEAREA 0.804 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585 1.62 2.515 1.79 ;
        RECT 0.585 1.165 0.915 1.62 ;
        RECT 1.845 1.35 2.515 1.62 ;
    END
    ANTENNAGATEAREA 0.804 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.99 0.255 4.175 0.425 ;
      RECT 3.84 0.425 4.175 0.5 ;
      RECT 1.97 0.67 3.16 0.84 ;
      RECT 2.99 0.425 3.16 0.67 ;
      RECT 1.97 0.35 2.3 0.67 ;
      RECT 2.495 2.905 3.675 3.075 ;
      RECT 3.395 2.36 3.675 2.905 ;
      RECT 3.395 2.19 4.685 2.36 ;
      RECT 4.345 2.36 4.685 2.98 ;
      RECT 1.545 2.47 1.795 2.98 ;
      RECT 1.545 2.3 2.825 2.47 ;
      RECT 2.495 2.47 2.825 2.905 ;
      RECT 2.685 1.35 3.125 1.68 ;
      RECT 0.245 1.96 2.855 2.13 ;
      RECT 2.685 1.68 2.855 1.96 ;
      RECT 0.245 0.84 0.415 1.96 ;
      RECT 1.065 2.13 1.315 2.98 ;
      RECT 0.245 0.67 1.22 0.84 ;
      RECT 0.89 0.35 1.22 0.67 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 3.845 2.53 4.175 3.245 ;
      RECT 1.995 2.64 2.325 3.245 ;
      RECT 0.115 2.3 0.445 3.245 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 0.115 0.085 0.71 0.5 ;
      RECT 1.39 0.085 1.72 0.84 ;
      RECT 2.48 0.085 2.82 0.5 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_xor2_2

MACRO scs8ls_xor2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985 2.285 6.315 2.455 ;
        RECT 2.985 2.455 3.315 2.735 ;
        RECT 3.885 2.455 4.215 2.735 ;
        RECT 2.985 2.19 3.315 2.285 ;
        RECT 6.145 2.12 6.315 2.285 ;
        RECT 6.145 1.95 8.505 2.12 ;
        RECT 8.335 1.18 8.505 1.95 ;
        RECT 4.105 1.01 8.505 1.18 ;
        RECT 4.105 0.85 4.275 1.01 ;
        RECT 6.835 0.595 7.165 1.01 ;
        RECT 7.845 0.595 8.015 1.01 ;
        RECT 3.21 0.68 4.275 0.85 ;
        RECT 3.21 0.47 3.54 0.68 ;
    END
    ANTENNADIFFAREA 1.5045 ;
  END X

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.805 1.55 8.165 1.78 ;
        RECT 5.805 1.78 5.975 1.945 ;
        RECT 5.885 1.35 8.165 1.55 ;
        RECT 2.03 1.945 5.975 2.02 ;
        RECT 3.485 2.02 5.975 2.115 ;
        RECT 2.03 1.85 3.655 1.945 ;
        RECT 2.03 1.47 2.36 1.85 ;
    END
    ANTENNAGATEAREA 1.638 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.52 5.635 1.775 ;
        RECT 3.765 1.35 5.635 1.52 ;
        RECT 3.765 1.19 3.935 1.35 ;
        RECT 2.87 1.02 3.935 1.19 ;
        RECT 2.87 0.77 3.04 1.02 ;
        RECT 1.275 0.75 3.04 0.77 ;
        RECT 0.515 0.6 3.04 0.75 ;
        RECT 0.515 0.75 0.685 1.42 ;
        RECT 0.515 0.58 1.445 0.6 ;
        RECT 0.44 1.42 1.11 1.75 ;
    END
    ANTENNAGATEAREA 1.638 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 6.405 0.255 8.525 0.425 ;
      RECT 8.195 0.425 8.525 0.84 ;
      RECT 4.445 0.67 6.655 0.84 ;
      RECT 6.405 0.425 6.655 0.67 ;
      RECT 4.445 0.35 4.695 0.67 ;
      RECT 5.385 0.35 5.715 0.67 ;
      RECT 7.335 0.425 7.665 0.84 ;
      RECT 1.11 2.905 2.34 3.075 ;
      RECT 2.01 2.19 2.34 2.905 ;
      RECT 1.11 2.09 1.36 2.905 ;
      RECT 0.16 1.92 1.36 2.09 ;
      RECT 0.16 2.09 0.49 2.98 ;
      RECT 4.415 2.625 6.655 2.795 ;
      RECT 6.485 2.795 6.655 2.98 ;
      RECT 6.485 2.46 6.655 2.625 ;
      RECT 6.485 2.29 8.535 2.46 ;
      RECT 7.305 2.46 7.635 2.98 ;
      RECT 8.205 2.46 8.535 2.98 ;
      RECT 2.535 2.19 2.785 2.905 ;
      RECT 3.515 2.625 3.685 2.905 ;
      RECT 2.535 2.905 4.665 3.075 ;
      RECT 4.415 2.795 4.665 2.905 ;
      RECT 5.375 2.795 5.705 2.98 ;
      RECT 2.53 1.36 3.595 1.68 ;
      RECT 0.855 1.19 1.105 1.25 ;
      RECT 1.56 1.19 1.81 2.735 ;
      RECT 0.855 0.92 1.105 0.94 ;
      RECT 2.53 1.19 2.7 1.36 ;
      RECT 0.855 0.94 2.7 1.19 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 5.89 2.965 6.22 3.245 ;
      RECT 6.855 2.63 7.105 3.245 ;
      RECT 7.835 2.63 8.005 3.245 ;
      RECT 0.69 2.26 0.94 3.245 ;
      RECT 4.855 2.965 5.185 3.245 ;
      RECT 0 -0.085 8.64 0.085 ;
      RECT 3.72 0.085 4.135 0.51 ;
      RECT 4.875 0.085 5.205 0.5 ;
      RECT 5.895 0.085 6.225 0.5 ;
      RECT 0.095 0.085 0.345 1.25 ;
      RECT 1.285 0.085 1.615 0.41 ;
      RECT 2.415 0.085 2.745 0.43 ;
    LAYER mcon ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
  END
END scs8ls_xor2_4

MACRO scs8ls_xor3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.755 0.4 9.005 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.96 1.18 1.285 1.75 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.875 1.18 7.205 1.685 ;
    END
    ANTENNAGATEAREA 0.381 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.92 1.35 5.25 1.78 ;
    END
    ANTENNAGATEAREA 0.693 ;
  END B

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 2.975 1.735 3.265 1.78 ;
      RECT 2.975 1.595 5.665 1.735 ;
      RECT 5.375 1.735 5.665 1.78 ;
      RECT 2.975 1.55 3.265 1.595 ;
      RECT 5.375 1.55 5.665 1.595 ;
      RECT 6.335 1.735 6.625 1.78 ;
      RECT 6.335 1.595 8.545 1.735 ;
      RECT 8.255 1.735 8.545 1.78 ;
      RECT 6.335 1.55 6.625 1.595 ;
      RECT 8.255 1.55 8.545 1.595 ;
    LAYER li1 ;
      RECT 6.025 2.905 7.605 3.075 ;
      RECT 7.435 2.525 7.605 2.905 ;
      RECT 7.435 2.195 7.985 2.525 ;
      RECT 7.815 0.86 7.985 2.195 ;
      RECT 7.815 0.4 8.065 0.86 ;
      RECT 6.025 1.82 6.195 2.905 ;
      RECT 5.805 1.53 6.195 1.82 ;
      RECT 3.725 1.435 4.055 1.735 ;
      RECT 3.725 0.765 3.895 1.435 ;
      RECT 3.725 0.595 4.805 0.765 ;
      RECT 4.58 0.765 4.805 1.13 ;
      RECT 4.58 1.13 4.75 2.98 ;
      RECT 5.775 0.255 7.645 0.425 ;
      RECT 7.475 0.425 7.645 1.855 ;
      RECT 6.875 1.855 7.645 2.025 ;
      RECT 6.875 2.025 7.205 2.735 ;
      RECT 3.385 0.255 5.145 0.425 ;
      RECT 4.975 0.425 5.145 0.85 ;
      RECT 4.975 0.85 6.025 1.02 ;
      RECT 5.775 0.425 6.025 0.85 ;
      RECT 1.93 2.565 3.555 2.735 ;
      RECT 1.93 1.94 2.26 2.565 ;
      RECT 3.385 0.425 3.555 2.565 ;
      RECT 6.365 1.55 6.705 2.735 ;
      RECT 6.535 0.935 6.705 1.55 ;
      RECT 2.965 1.875 3.215 2.395 ;
      RECT 3.02 0.46 3.215 1.875 ;
      RECT 2.135 0.29 3.215 0.46 ;
      RECT 2.135 0.46 2.385 1.09 ;
      RECT 8.255 1.35 8.585 1.78 ;
      RECT 6.195 0.595 7.305 0.765 ;
      RECT 6.885 0.765 7.305 0.925 ;
      RECT 5.405 1.99 5.855 2.84 ;
      RECT 5.405 1.95 5.625 1.99 ;
      RECT 5.42 1.36 5.625 1.95 ;
      RECT 5.42 1.19 6.365 1.36 ;
      RECT 6.195 0.765 6.365 1.19 ;
      RECT 1.37 2.905 3.895 3.075 ;
      RECT 3.725 2.755 3.895 2.905 ;
      RECT 1.37 2.09 1.7 2.905 ;
      RECT 3.725 1.905 4.395 2.755 ;
      RECT 0.425 1.94 1.7 2.09 ;
      RECT 4.225 1.265 4.395 1.905 ;
      RECT 0.425 1.92 1.625 1.94 ;
      RECT 4.065 0.935 4.395 1.265 ;
      RECT 1.455 1 1.625 1.92 ;
      RECT 0.425 1.47 0.75 1.92 ;
      RECT 0.085 0.66 1.965 0.83 ;
      RECT 1.795 0.83 1.965 1.26 ;
      RECT 1.795 1.26 2.76 1.43 ;
      RECT 2.43 1.43 2.76 2.395 ;
      RECT 2.59 1.09 2.76 1.26 ;
      RECT 2.59 0.63 2.85 1.09 ;
      RECT 0.085 2.26 0.6 2.98 ;
      RECT 0.085 1.3 0.255 2.26 ;
      RECT 0.085 0.83 0.445 1.3 ;
      RECT 0.085 0.65 0.445 0.66 ;
      RECT 0 3.245 9.12 3.415 ;
      RECT 0.77 2.26 1.1 3.245 ;
      RECT 4.95 1.95 5.2 3.245 ;
      RECT 8.225 1.95 8.555 3.245 ;
      RECT 0 -0.085 9.12 0.085 ;
      RECT 0.625 0.085 1.195 0.49 ;
      RECT 5.315 0.085 5.565 0.68 ;
      RECT 8.245 0.085 8.575 1.18 ;
    LAYER mcon ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.395 1.58 6.565 1.75 ;
      RECT 5.435 1.58 5.605 1.75 ;
      RECT 3.035 1.58 3.205 1.75 ;
      RECT 8.315 1.58 8.485 1.75 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
  END
END scs8ls_xor3_1

MACRO scs8ls_xor3_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.705 0.37 9.035 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955 1.18 1.285 1.75 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.875 1.18 7.125 1.685 ;
    END
    ANTENNAGATEAREA 0.381 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.92 1.18 5.25 1.55 ;
    END
    ANTENNAGATEAREA 0.693 ;
  END B

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 6.335 2.105 6.625 2.15 ;
      RECT 6.335 1.965 8.545 2.105 ;
      RECT 8.255 2.105 8.545 2.15 ;
      RECT 6.335 1.92 6.625 1.965 ;
      RECT 8.255 1.92 8.545 1.965 ;
      RECT 2.975 2.105 3.265 2.15 ;
      RECT 2.975 1.965 5.665 2.105 ;
      RECT 5.375 2.105 5.665 2.15 ;
      RECT 2.975 1.92 3.265 1.965 ;
      RECT 5.375 1.92 5.665 1.965 ;
    LAYER li1 ;
      RECT 8.315 1.65 8.525 2.15 ;
      RECT 8.195 1.32 8.525 1.65 ;
      RECT 3.725 1.435 4.055 1.735 ;
      RECT 3.725 0.765 3.895 1.435 ;
      RECT 3.725 0.595 4.805 0.765 ;
      RECT 4.58 0.765 4.805 1.01 ;
      RECT 4.58 1.01 4.75 2.98 ;
      RECT 6.01 2.905 7.45 3.075 ;
      RECT 7.28 2.5 7.45 2.905 ;
      RECT 7.28 2.195 7.805 2.5 ;
      RECT 7.635 1.605 7.805 2.195 ;
      RECT 7.635 1.435 8.025 1.605 ;
      RECT 7.775 0.37 8.025 1.435 ;
      RECT 6.01 1.685 6.18 2.905 ;
      RECT 5.85 1.355 6.18 1.685 ;
      RECT 5.775 0.255 7.605 0.425 ;
      RECT 7.435 0.425 7.605 1.095 ;
      RECT 7.295 1.095 7.605 1.265 ;
      RECT 7.295 1.265 7.465 1.855 ;
      RECT 6.785 1.855 7.465 2.025 ;
      RECT 6.785 2.025 7.05 2.69 ;
      RECT 3.385 0.255 5.145 0.425 ;
      RECT 4.975 0.425 5.145 0.675 ;
      RECT 4.975 0.675 6.025 0.845 ;
      RECT 5.775 0.425 6.025 0.675 ;
      RECT 1.85 2.565 3.555 2.735 ;
      RECT 1.85 2.075 2.18 2.565 ;
      RECT 3.385 0.425 3.555 2.565 ;
      RECT 6.35 1.525 6.6 2.7 ;
      RECT 6.35 1.355 6.705 1.525 ;
      RECT 6.535 0.935 6.705 1.355 ;
      RECT 2.885 1.875 3.215 2.395 ;
      RECT 3.045 0.595 3.215 1.875 ;
      RECT 2.135 0.425 3.215 0.595 ;
      RECT 2.135 0.595 2.305 1.225 ;
      RECT 6.195 0.595 7.265 0.765 ;
      RECT 6.885 0.765 7.265 0.925 ;
      RECT 5.405 1.92 5.84 2.98 ;
      RECT 5.51 1.185 5.68 1.92 ;
      RECT 5.51 1.015 6.365 1.185 ;
      RECT 6.195 0.765 6.365 1.015 ;
      RECT 0.085 0.66 1.965 0.83 ;
      RECT 1.795 0.83 1.965 1.395 ;
      RECT 1.795 1.395 2.68 1.565 ;
      RECT 2.35 1.565 2.68 2.395 ;
      RECT 2.51 1.225 2.68 1.395 ;
      RECT 2.51 0.765 2.875 1.225 ;
      RECT 0.085 2.26 0.595 2.955 ;
      RECT 0.085 1.275 0.255 2.26 ;
      RECT 0.085 0.83 0.445 1.275 ;
      RECT 0.085 0.65 0.445 0.66 ;
      RECT 1.31 2.905 3.895 3.075 ;
      RECT 3.725 2.755 3.895 2.905 ;
      RECT 1.31 2.09 1.64 2.905 ;
      RECT 3.725 1.905 4.395 2.755 ;
      RECT 0.425 2.075 1.64 2.09 ;
      RECT 4.225 1.265 4.395 1.905 ;
      RECT 0.425 1.92 1.625 2.075 ;
      RECT 4.065 0.935 4.395 1.265 ;
      RECT 1.455 1 1.625 1.92 ;
      RECT 0.425 1.445 0.745 1.92 ;
      RECT 0 3.245 9.6 3.415 ;
      RECT 9.235 1.82 9.485 3.245 ;
      RECT 7.975 2.32 8.53 3.245 ;
      RECT 0.765 2.26 1.095 3.245 ;
      RECT 4.95 1.82 5.2 3.245 ;
      RECT 7.975 1.82 8.145 2.32 ;
      RECT 0 -0.085 9.6 0.085 ;
      RECT 9.215 0.085 9.465 1.15 ;
      RECT 0.625 0.085 1.195 0.49 ;
      RECT 5.315 0.085 5.565 0.505 ;
      RECT 8.205 0.085 8.535 1.15 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.395 1.95 6.565 2.12 ;
      RECT 5.435 1.95 5.605 2.12 ;
      RECT 8.315 1.95 8.485 2.12 ;
      RECT 3.035 1.95 3.205 2.12 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
  END
END scs8ls_xor3_2

MACRO scs8ls_xor3_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.91 1.18 1.285 1.67 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.81 1.45 7.07 1.78 ;
    END
    ANTENNAGATEAREA 0.381 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.91 1.18 5.24 1.55 ;
    END
    ANTENNAGATEAREA 0.693 ;
  END B

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.665 1.55 9.995 2.98 ;
        RECT 9.665 1.47 9.94 1.55 ;
        RECT 8.955 1.3 9.94 1.47 ;
        RECT 8.955 1.47 9.125 1.82 ;
        RECT 8.955 1.085 9.16 1.3 ;
        RECT 9.69 0.35 9.94 1.3 ;
        RECT 8.685 1.82 9.125 2.98 ;
        RECT 8.83 0.35 9.16 1.085 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 6.335 2.105 6.625 2.15 ;
      RECT 6.335 1.965 8.545 2.105 ;
      RECT 8.255 2.105 8.545 2.15 ;
      RECT 6.335 1.92 6.625 1.965 ;
      RECT 8.255 1.92 8.545 1.965 ;
      RECT 2.495 2.105 2.785 2.15 ;
      RECT 2.495 1.965 5.665 2.105 ;
      RECT 5.375 2.105 5.665 2.15 ;
      RECT 2.495 1.92 2.785 1.965 ;
      RECT 5.375 1.92 5.665 1.965 ;
    LAYER li1 ;
      RECT 0 -0.085 10.56 0.085 ;
      RECT 10.12 0.085 10.45 1.13 ;
      RECT 0.625 0.085 1.035 0.41 ;
      RECT 5.25 0.085 5.5 0.61 ;
      RECT 8.33 0.085 8.66 1.085 ;
      RECT 9.34 0.085 9.51 1.13 ;
      RECT 0 3.245 10.56 3.415 ;
      RECT 10.195 1.82 10.445 3.245 ;
      RECT 7.945 2.33 8.5 3.245 ;
      RECT 0.565 2.18 0.895 3.245 ;
      RECT 4.905 1.82 5.235 3.245 ;
      RECT 7.945 1.82 8.115 2.33 ;
      RECT 9.295 1.82 9.465 3.245 ;
      RECT 7.92 1.255 8.785 1.585 ;
      RECT 8.285 1.585 8.515 2.15 ;
      RECT 5.965 2.905 7.5 3.075 ;
      RECT 7.33 2.71 7.5 2.905 ;
      RECT 7.33 2.29 7.75 2.71 ;
      RECT 7.58 0.745 7.75 2.29 ;
      RECT 7.58 0.415 8.15 0.745 ;
      RECT 5.965 1.75 6.135 2.905 ;
      RECT 5.775 1.46 6.135 1.75 ;
      RECT 5.71 0.255 7.41 0.425 ;
      RECT 7.24 0.425 7.41 1.95 ;
      RECT 6.835 1.95 7.41 2.12 ;
      RECT 6.835 2.12 7.085 2.735 ;
      RECT 3.315 0.255 5.08 0.425 ;
      RECT 4.91 0.425 5.08 0.78 ;
      RECT 4.91 0.78 5.96 0.95 ;
      RECT 5.71 0.425 5.96 0.78 ;
      RECT 1.6 2.565 3.485 2.735 ;
      RECT 1.6 2.18 1.93 2.565 ;
      RECT 3.315 0.425 3.485 2.565 ;
      RECT 6.13 0.595 7.07 0.765 ;
      RECT 6.82 0.765 7.07 1.275 ;
      RECT 5.405 1.92 5.795 2.8 ;
      RECT 5.435 1.29 5.605 1.92 ;
      RECT 5.435 1.12 6.3 1.29 ;
      RECT 6.13 0.765 6.3 1.12 ;
      RECT 6.305 1.92 6.64 2.735 ;
      RECT 6.47 0.935 6.64 1.92 ;
      RECT 3.655 1.435 3.985 1.735 ;
      RECT 3.655 0.765 3.825 1.435 ;
      RECT 3.655 0.595 4.74 0.765 ;
      RECT 4.535 0.765 4.74 1.13 ;
      RECT 4.535 1.13 4.705 2.98 ;
      RECT 1.065 2.905 3.825 3.075 ;
      RECT 3.655 2.755 3.825 2.905 ;
      RECT 1.065 2.01 1.395 2.905 ;
      RECT 3.655 1.905 4.325 2.755 ;
      RECT 0.425 1.84 1.625 2.01 ;
      RECT 4.155 1.265 4.325 1.905 ;
      RECT 1.455 0.92 1.625 1.84 ;
      RECT 3.995 0.935 4.325 1.265 ;
      RECT 0.425 1.47 0.7 1.84 ;
      RECT 2.555 1.875 3.145 2.395 ;
      RECT 2.975 0.62 3.145 1.875 ;
      RECT 2.135 0.45 3.145 0.62 ;
      RECT 2.135 0.62 2.385 1.25 ;
      RECT 0.085 0.58 1.965 0.75 ;
      RECT 1.795 0.75 1.965 1.42 ;
      RECT 1.795 1.42 2.805 1.59 ;
      RECT 2.135 1.59 2.385 2.395 ;
      RECT 2.555 0.79 2.805 1.42 ;
      RECT 0.085 2.18 0.365 2.98 ;
      RECT 0.085 1.25 0.255 2.18 ;
      RECT 0.085 0.75 0.445 1.25 ;
      RECT 0.085 0.57 0.445 0.58 ;
    LAYER mcon ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 1.95 8.485 2.12 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 1.95 6.565 2.12 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 1.95 5.605 2.12 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 1.95 2.725 2.12 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_xor3_4

MACRO scs8ls_or4bb_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.345 0.35 4.715 1.13 ;
        RECT 4.545 1.13 4.715 1.82 ;
        RECT 4.24 1.82 4.715 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.35 3.835 1.78 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.965 1.35 3.295 2.89 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END B

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.3 0.455 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END CN

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.05 1.315 1.72 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END DN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 3.74 1.95 4.07 3.245 ;
      RECT 0.615 2.65 0.945 3.245 ;
      RECT 0.115 2.31 1.285 2.48 ;
      RECT 1.115 2.48 1.285 2.905 ;
      RECT 1.115 2.905 2.755 3.075 ;
      RECT 2.425 1.19 2.755 2.905 ;
      RECT 0.115 2.48 0.445 2.98 ;
      RECT 0.115 2.1 0.795 2.31 ;
      RECT 0.625 1.13 0.795 2.1 ;
      RECT 0.14 0.96 0.795 1.13 ;
      RECT 0.14 0.35 0.47 0.96 ;
      RECT 4.005 1.3 4.375 1.63 ;
      RECT 2.075 1.01 4.175 1.02 ;
      RECT 3.31 1.02 4.175 1.18 ;
      RECT 2.075 0.85 3.64 1.01 ;
      RECT 4.005 1.18 4.175 1.3 ;
      RECT 3.31 0.35 3.64 0.85 ;
      RECT 1.845 1.87 2.245 2.735 ;
      RECT 2.075 1.02 2.245 1.87 ;
      RECT 2.245 0.35 2.575 0.85 ;
      RECT 1.15 1.89 1.655 2.14 ;
      RECT 1.485 1.7 1.655 1.89 ;
      RECT 1.485 1.03 1.905 1.7 ;
      RECT 1.485 0.88 1.655 1.03 ;
      RECT 1.14 0.35 1.655 0.88 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 0.64 0.085 0.97 0.79 ;
      RECT 1.825 0.085 2.075 0.68 ;
      RECT 2.745 0.085 3.14 0.68 ;
      RECT 3.81 0.085 4.14 0.84 ;
    LAYER mcon ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_or4bb_1

MACRO scs8ls_or4bb_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.47 3.925 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.15 0.255 3.715 0.57 ;
        RECT 3.485 0.57 3.715 0.67 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.435 1.3 4.695 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END CN

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 0.55 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END DN

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.06 0.44 1.315 1.18 ;
        RECT 1.06 1.18 1.23 1.85 ;
        RECT 1.06 1.85 1.39 2.1 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 0.605 2.61 0.935 3.245 ;
      RECT 1.51 2.61 1.84 3.245 ;
      RECT 3.82 2.31 4.15 3.245 ;
      RECT 1.56 1.13 3.735 1.3 ;
      RECT 3.405 0.84 3.735 1.13 ;
      RECT 2.05 2.78 2.38 2.98 ;
      RECT 2.05 2.61 2.605 2.78 ;
      RECT 2.435 1.3 2.605 2.61 ;
      RECT 1.56 1.3 1.73 1.35 ;
      RECT 2.31 0.58 2.64 1.13 ;
      RECT 1.4 1.35 1.73 1.68 ;
      RECT 0.105 2.27 2.265 2.44 ;
      RECT 1.97 1.47 2.265 2.27 ;
      RECT 0.105 2.44 0.435 2.98 ;
      RECT 0.105 2.1 0.89 2.27 ;
      RECT 0.72 1.18 0.89 2.1 ;
      RECT 0.12 1.01 0.89 1.18 ;
      RECT 0.12 0.67 0.45 1.01 ;
      RECT 4.36 2.14 4.69 2.82 ;
      RECT 2.775 1.97 4.69 2.14 ;
      RECT 4.095 1.95 4.69 1.97 ;
      RECT 4.095 0.96 4.685 1.13 ;
      RECT 4.435 0.435 4.685 0.96 ;
      RECT 4.095 1.13 4.265 1.95 ;
      RECT 2.775 1.47 3.07 1.97 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 3.925 0.085 4.255 0.79 ;
      RECT 2.81 0.085 2.98 0.74 ;
      RECT 1.575 0.085 2.035 0.91 ;
      RECT 2.81 0.74 3.195 0.96 ;
      RECT 0.63 0.085 0.88 0.84 ;
    LAYER mcon ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_or4bb_2

MACRO scs8ls_or4bb_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.45 7.075 1.78 ;
    END
    ANTENNAGATEAREA 0.411 ;
  END B

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.18 1.45 2.05 ;
        RECT 1.085 2.05 2.525 2.22 ;
        RECT 1.12 0.75 1.45 1.18 ;
        RECT 1.12 0.58 2.775 0.75 ;
        RECT 2.14 0.42 2.775 0.58 ;
        RECT 1.12 0.35 1.45 0.58 ;
    END
    ANTENNADIFFAREA 1.6775 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.525 1.18 8.535 1.55 ;
    END
    ANTENNAGATEAREA 0.411 ;
  END A

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.375 1.35 3.715 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END CN

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.35 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END DN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 7.245 1.95 8.525 2.24 ;
      RECT 7.245 2.24 7.575 2.905 ;
      RECT 8.195 1.94 8.525 1.95 ;
      RECT 6.345 2.905 7.575 3.075 ;
      RECT 6.345 2.44 6.675 2.905 ;
      RECT 8.25 2.24 8.525 2.99 ;
      RECT 4.835 2.98 6.115 3.075 ;
      RECT 3.935 2.905 6.115 2.98 ;
      RECT 3.935 2.63 5.165 2.905 ;
      RECT 5.865 2.44 6.115 2.905 ;
      RECT 5.335 2.27 5.665 2.735 ;
      RECT 5.335 2.1 7.045 2.27 ;
      RECT 6.875 2.27 7.045 2.735 ;
      RECT 6.575 1.95 7.045 2.1 ;
      RECT 1.62 0.92 4.275 1.09 ;
      RECT 3.945 1.09 4.275 1.25 ;
      RECT 0.085 2.39 2.865 2.56 ;
      RECT 2.695 1.88 2.865 2.39 ;
      RECT 1.62 1.71 2.865 1.88 ;
      RECT 0.085 2.56 0.445 2.86 ;
      RECT 0.085 1.95 0.445 2.39 ;
      RECT 0.085 0.45 0.445 1.13 ;
      RECT 0.085 1.13 0.255 1.95 ;
      RECT 1.62 1.09 1.79 1.71 ;
      RECT 5.975 1.09 7.355 1.26 ;
      RECT 7.025 0.35 7.355 1.09 ;
      RECT 3.035 2.29 4.715 2.46 ;
      RECT 4.385 1.93 4.715 2.29 ;
      RECT 4.385 1.76 6.145 1.93 ;
      RECT 5.975 1.26 6.145 1.76 ;
      RECT 4.785 0.35 6.28 1.09 ;
      RECT 3.035 1.54 3.205 2.29 ;
      RECT 1.96 1.26 3.205 1.54 ;
      RECT 3.375 1.95 4.055 2.12 ;
      RECT 3.885 1.59 4.055 1.95 ;
      RECT 3.885 1.42 5.805 1.59 ;
      RECT 4.445 1.26 5.805 1.42 ;
      RECT 4.445 0.75 4.615 1.26 ;
      RECT 3.455 0.58 4.615 0.75 ;
      RECT 3.455 0.45 3.785 0.58 ;
      RECT 0 -0.085 8.64 0.085 ;
      RECT 2.945 0.085 3.275 0.75 ;
      RECT 4.015 0.085 4.605 0.41 ;
      RECT 6.45 0.085 6.78 0.92 ;
      RECT 7.64 0.085 8.31 0.985 ;
      RECT 0.615 0.085 0.915 1.13 ;
      RECT 1.63 0.085 1.96 0.41 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 0.65 2.73 0.995 3.245 ;
      RECT 1.565 2.73 1.99 3.245 ;
      RECT 2.84 2.73 3.17 3.245 ;
      RECT 7.745 2.41 8.075 3.245 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
  END
END scs8ls_or4bb_4

MACRO scs8ls_sdfbbn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 16.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.355 1.82 16.715 2.98 ;
        RECT 16.545 1.05 16.715 1.82 ;
        RECT 16.335 0.35 16.715 1.05 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END Q

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.075 1.19 14.38 1.55 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END RESETB

  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.47 1.35 3.8 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLKN

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.89 1.82 15.275 2.98 ;
        RECT 15.105 1.13 15.275 1.82 ;
        RECT 14.915 0.35 15.275 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END QN

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.205 0.55 1.875 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805 1.205 1.315 1.875 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.48 1.815 1.81 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 16.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 16.8 3.575 ;
    END
  END vpwr

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 8.255 1.965 11.905 2.105 ;
        RECT 11.615 2.105 11.905 2.15 ;
        RECT 11.615 1.92 11.905 1.965 ;
        RECT 8.255 2.105 8.545 2.15 ;
        RECT 8.255 1.92 8.545 1.965 ;
    END
    ANTENNAGATEAREA 0.4695 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.541 LAYER met1 ;
  END SETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 12.465 0.79 13.565 0.96 ;
      RECT 12.465 0.595 12.795 0.79 ;
      RECT 15.45 1.22 16.375 1.55 ;
      RECT 15.45 1.55 15.7 2.78 ;
      RECT 15.45 0.35 15.725 1.22 ;
      RECT 11.63 1.47 11.96 2.12 ;
      RECT 0 3.245 16.8 3.415 ;
      RECT 15.905 1.9 16.155 3.245 ;
      RECT 10.9 2.97 11.23 3.245 ;
      RECT 11.995 2.97 12.325 3.245 ;
      RECT 8.125 2.65 8.295 3.245 ;
      RECT 14 2.55 14.69 3.245 ;
      RECT 9.05 2.47 9.38 3.245 ;
      RECT 5.02 2.465 5.27 3.245 ;
      RECT 0.565 2.385 0.895 3.245 ;
      RECT 2.47 2.3 2.72 3.245 ;
      RECT 3.93 2.29 4.18 3.245 ;
      RECT 0 -0.085 16.8 0.085 ;
      RECT 15.905 0.085 16.155 1.05 ;
      RECT 0.14 0.085 0.47 1.035 ;
      RECT 1.89 0.085 2.22 0.97 ;
      RECT 3.8 0.085 4.13 0.41 ;
      RECT 5.3 0.085 5.63 1.035 ;
      RECT 8.795 0.085 9.125 1.08 ;
      RECT 11.415 0.085 11.755 0.41 ;
      RECT 14.415 0.085 14.735 0.68 ;
      RECT 8.285 1.96 8.49 2.14 ;
      RECT 8.285 1.79 8.99 1.96 ;
      RECT 8.66 1.63 8.99 1.79 ;
      RECT 9.725 1.555 10.07 1.94 ;
      RECT 9.725 1.26 11 1.555 ;
      RECT 11.935 0.425 12.265 0.96 ;
      RECT 11.935 0.255 13.225 0.425 ;
      RECT 12.975 0.425 13.225 0.62 ;
      RECT 13.61 1.79 14.13 2.04 ;
      RECT 13.61 1.3 13.78 1.79 ;
      RECT 11.51 1.13 13.905 1.3 ;
      RECT 12.2 1.3 12.53 1.55 ;
      RECT 11.51 0.75 11.68 1.13 ;
      RECT 13.735 0.67 13.905 1.13 ;
      RECT 10.75 0.58 11.68 0.75 ;
      RECT 10.75 0.535 10.92 0.58 ;
      RECT 9.385 0.365 10.92 0.535 ;
      RECT 9.385 0.535 9.555 1.29 ;
      RECT 8.1 1.29 9.555 1.46 ;
      RECT 8.1 1.46 8.43 1.62 ;
      RECT 4.38 1.84 4.78 2.98 ;
      RECT 4.61 1.72 4.78 1.84 ;
      RECT 4.61 1.55 6.71 1.72 ;
      RECT 5.405 1.72 6.71 1.8 ;
      RECT 6.38 1.47 6.71 1.55 ;
      RECT 4.61 1.17 4.79 1.55 ;
      RECT 5.405 1.8 5.755 1.905 ;
      RECT 4.31 0.92 4.79 1.17 ;
      RECT 6.365 2.48 6.695 2.735 ;
      RECT 6.365 2.31 7.59 2.48 ;
      RECT 7.42 0.96 7.59 2.31 ;
      RECT 6.595 0.79 7.59 0.96 ;
      RECT 6.595 0.425 6.925 0.79 ;
      RECT 5.8 0.255 6.925 0.425 ;
      RECT 5.8 0.425 5.97 1.205 ;
      RECT 4.96 1.205 5.97 1.375 ;
      RECT 4.96 0.75 5.13 1.205 ;
      RECT 3.23 0.58 5.13 0.75 ;
      RECT 3.23 0.425 3.4 0.58 ;
      RECT 2.39 0.255 3.4 0.425 ;
      RECT 2.39 0.425 2.56 1.14 ;
      RECT 1.485 1.14 2.56 1.31 ;
      RECT 1.985 1.31 2.155 1.98 ;
      RECT 1.485 1.035 1.655 1.14 ;
      RECT 1.545 1.98 2.155 2.15 ;
      RECT 0.96 0.865 1.655 1.035 ;
      RECT 1.545 2.15 1.715 2.3 ;
      RECT 1.465 2.3 1.715 2.735 ;
      RECT 0.96 0.575 1.29 0.865 ;
      RECT 7.15 0.425 7.48 0.62 ;
      RECT 7.15 0.255 8.59 0.425 ;
      RECT 8.26 0.425 8.59 1.08 ;
      RECT 1.065 2.905 2.245 3.075 ;
      RECT 1.915 2.32 2.245 2.905 ;
      RECT 1.065 2.215 1.235 2.905 ;
      RECT 0.115 2.045 1.235 2.215 ;
      RECT 0.115 2.215 0.395 2.98 ;
      RECT 3.48 2.12 3.73 2.98 ;
      RECT 3.48 1.95 4.14 2.12 ;
      RECT 3.97 1.67 4.14 1.95 ;
      RECT 3.97 1.34 4.44 1.67 ;
      RECT 3.97 1.17 4.14 1.34 ;
      RECT 3.29 0.92 4.14 1.17 ;
      RECT 2.89 2.3 3.25 2.98 ;
      RECT 2.89 1.81 3.06 2.3 ;
      RECT 2.51 1.48 3.06 1.81 ;
      RECT 2.73 0.595 3.06 1.48 ;
      RECT 5.865 2.245 6.195 2.735 ;
      RECT 6.025 2.14 6.195 2.245 ;
      RECT 6.025 1.97 7.25 2.14 ;
      RECT 6.92 1.3 7.25 1.97 ;
      RECT 6.17 1.13 7.25 1.3 ;
      RECT 6.17 0.595 6.42 1.13 ;
      RECT 5.44 2.905 7.505 3.075 ;
      RECT 6.925 2.82 7.505 2.905 ;
      RECT 5.44 2.295 5.61 2.905 ;
      RECT 6.925 2.65 7.93 2.82 ;
      RECT 4.95 2.125 5.61 2.295 ;
      RECT 7.76 2.48 7.93 2.65 ;
      RECT 4.95 1.965 5.215 2.125 ;
      RECT 7.76 2.31 8.83 2.48 ;
      RECT 8.495 2.48 8.83 2.98 ;
      RECT 8.66 2.3 8.83 2.31 ;
      RECT 7.76 1.08 7.93 2.31 ;
      RECT 8.66 2.13 9.53 2.3 ;
      RECT 7.76 0.595 8.09 1.08 ;
      RECT 9.2 1.63 9.53 2.13 ;
      RECT 9.89 2.28 10.22 2.98 ;
      RECT 9.89 2.11 10.41 2.28 ;
      RECT 10.24 1.895 10.41 2.11 ;
      RECT 10.24 1.725 11.34 1.895 ;
      RECT 11.17 1.895 11.34 2.29 ;
      RECT 11.17 1.09 11.34 1.725 ;
      RECT 11.17 2.29 12.78 2.46 ;
      RECT 9.745 0.92 11.34 1.09 ;
      RECT 12.61 1.89 12.78 2.29 ;
      RECT 9.745 0.705 10.58 0.92 ;
      RECT 12.61 1.72 13.44 1.89 ;
      RECT 12.77 1.47 13.44 1.72 ;
      RECT 14.55 1.3 14.935 1.63 ;
      RECT 12.95 2.21 14.72 2.38 ;
      RECT 14.55 1.63 14.72 2.21 ;
      RECT 14.55 1.02 14.72 1.3 ;
      RECT 14.075 0.85 14.72 1.02 ;
      RECT 14.075 0.5 14.245 0.85 ;
      RECT 13.395 0.33 14.245 0.5 ;
      RECT 11.46 2.8 11.79 2.98 ;
      RECT 10.665 2.63 13.28 2.8 ;
      RECT 12.95 2.8 13.28 2.98 ;
      RECT 12.95 2.38 13.28 2.63 ;
      RECT 10.665 2.065 10.995 2.63 ;
      RECT 12.95 2.06 13.28 2.21 ;
      RECT 13.395 0.5 13.565 0.79 ;
    LAYER mcon ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.315 1.95 8.485 2.12 ;
      RECT 5.435 1.58 5.605 1.75 ;
      RECT 9.755 1.58 9.925 1.75 ;
      RECT 11.675 1.95 11.845 2.12 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 14.555 -0.085 14.725 0.085 ;
    LAYER met1 ;
      RECT 5.375 1.735 5.665 1.78 ;
      RECT 5.375 1.595 9.985 1.735 ;
      RECT 9.695 1.735 9.985 1.78 ;
      RECT 5.375 1.55 5.665 1.595 ;
      RECT 9.695 1.55 9.985 1.595 ;
  END
END scs8ls_sdfbbn_1

MACRO scs8ls_sdfbbn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 18.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.945 1.505 14.275 1.835 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END RESETB

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 17.395 1.82 17.705 2.98 ;
        RECT 17.535 1.05 17.705 1.82 ;
        RECT 17.37 0.35 17.705 1.05 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.375 1.55 15.715 1.78 ;
        RECT 15.375 1.78 15.625 2.98 ;
        RECT 15.375 1.22 15.61 1.55 ;
        RECT 15.28 0.35 15.61 1.22 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END QN

  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.35 3.895 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLKN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.46 1.815 1.79 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805 1.125 1.315 1.795 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.125 0.55 2.135 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 18.24 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 18.24 3.575 ;
    END
  END vpwr

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 9.215 1.595 12.385 1.735 ;
        RECT 12.095 1.735 12.385 1.78 ;
        RECT 12.095 1.55 12.385 1.595 ;
        RECT 9.215 1.735 9.505 1.78 ;
        RECT 9.215 1.55 9.505 1.595 ;
    END
    ANTENNAGATEAREA 0.4695 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.205 LAYER met1 ;
  END SETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 14.485 1.005 14.655 1.43 ;
      RECT 14.32 0.835 14.655 1.005 ;
      RECT 12.835 0.665 14.49 0.835 ;
      RECT 13.185 2.675 13.435 2.98 ;
      RECT 13.185 2.43 13.435 2.505 ;
      RECT 11.08 2.26 13.435 2.43 ;
      RECT 11.805 2.43 12.135 2.98 ;
      RECT 11.08 2.09 11.41 2.26 ;
      RECT 13.185 2.06 13.435 2.26 ;
      RECT 12.835 0.835 13.085 0.96 ;
      RECT 12.835 0.595 13.085 0.665 ;
      RECT 16.34 1.55 16.7 2.94 ;
      RECT 16.34 1.22 17.365 1.55 ;
      RECT 16.34 0.54 16.67 1.22 ;
      RECT 4.405 1.84 4.785 2.98 ;
      RECT 4.615 1.35 4.785 1.84 ;
      RECT 4.615 1.18 6.115 1.35 ;
      RECT 5.595 1.35 6.115 1.525 ;
      RECT 4.69 0.595 4.94 1.18 ;
      RECT 5.595 1.525 6.825 1.84 ;
      RECT 6.495 1.84 6.825 1.855 ;
      RECT 11.955 1.18 12.325 1.75 ;
      RECT 0 -0.085 18.24 0.085 ;
      RECT 17.88 0.085 18.13 1.13 ;
      RECT 15.78 0.085 16.11 1.13 ;
      RECT 16.87 0.085 17.2 1.05 ;
      RECT 2.18 0.085 2.43 0.95 ;
      RECT 3.93 0.085 4.18 0.49 ;
      RECT 5.45 0.085 5.72 0.67 ;
      RECT 9.055 0.085 9.385 0.94 ;
      RECT 11.68 0.085 12.055 0.43 ;
      RECT 14.825 0.085 15.11 1.13 ;
      RECT 0.14 0.085 0.47 0.955 ;
      RECT 0 3.245 18.24 3.415 ;
      RECT 17.875 1.82 18.125 3.245 ;
      RECT 15.825 1.95 16.155 3.245 ;
      RECT 16.895 1.82 17.225 3.245 ;
      RECT 14.28 2.845 15.17 3.245 ;
      RECT 14.825 1.95 15.17 2.845 ;
      RECT 0.565 2.645 0.895 3.245 ;
      RECT 11.23 2.6 11.56 3.245 ;
      RECT 12.305 2.6 12.635 3.245 ;
      RECT 8.365 2.465 8.695 3.245 ;
      RECT 4.965 2.35 5.215 3.245 ;
      RECT 2.415 2.3 2.745 3.245 ;
      RECT 3.875 2.29 4.205 3.245 ;
      RECT 9.465 2.29 9.795 3.245 ;
      RECT 8.79 1.45 9.445 1.78 ;
      RECT 12.235 0.425 12.655 0.6 ;
      RECT 12.235 0.255 13.595 0.425 ;
      RECT 13.265 0.425 13.595 0.495 ;
      RECT 10.155 1.58 10.485 1.755 ;
      RECT 10.155 1.28 11.385 1.58 ;
      RECT 10.155 1.18 10.485 1.28 ;
      RECT 13.605 2.005 14.075 2.335 ;
      RECT 13.605 1.3 14.15 1.335 ;
      RECT 12.495 1.13 14.15 1.3 ;
      RECT 13.605 1.005 14.15 1.13 ;
      RECT 13.605 1.335 13.775 2.005 ;
      RECT 12.495 1.3 12.825 1.55 ;
      RECT 12.495 0.94 12.665 1.13 ;
      RECT 11.895 0.77 12.665 0.94 ;
      RECT 11.34 0.6 12.065 0.77 ;
      RECT 11.34 0.43 11.51 0.6 ;
      RECT 9.555 0.26 11.51 0.43 ;
      RECT 9.555 0.43 9.725 1.11 ;
      RECT 8.45 1.11 9.725 1.28 ;
      RECT 8.45 1.28 8.62 1.285 ;
      RECT 8.215 1.285 8.62 1.955 ;
      RECT 8.45 0.605 8.885 0.935 ;
      RECT 8.45 0.435 8.62 0.605 ;
      RECT 7.345 0.265 8.62 0.435 ;
      RECT 7.345 0.435 7.77 0.675 ;
      RECT 5.84 2.21 6.17 2.735 ;
      RECT 5.84 2.04 7.365 2.21 ;
      RECT 7.035 1.355 7.365 2.04 ;
      RECT 6.285 1.185 7.365 1.355 ;
      RECT 6.285 0.605 6.615 1.185 ;
      RECT 6.34 2.55 6.67 2.735 ;
      RECT 6.34 2.38 7.705 2.55 ;
      RECT 7.535 1.015 7.705 2.38 ;
      RECT 6.785 0.845 7.705 1.015 ;
      RECT 6.785 0.435 7.115 0.845 ;
      RECT 5.945 0.265 7.115 0.435 ;
      RECT 5.945 0.435 6.115 0.84 ;
      RECT 5.11 0.84 6.115 1.01 ;
      RECT 5.11 0.425 5.28 0.84 ;
      RECT 4.35 0.255 5.28 0.425 ;
      RECT 4.35 0.425 4.52 0.66 ;
      RECT 3.365 0.66 4.52 0.83 ;
      RECT 3.365 0.425 3.535 0.66 ;
      RECT 2.6 0.255 3.535 0.425 ;
      RECT 2.6 0.425 2.77 1.12 ;
      RECT 1.485 1.12 2.77 1.29 ;
      RECT 1.985 1.29 2.155 1.96 ;
      RECT 1.485 0.955 1.69 1.12 ;
      RECT 1.485 1.96 2.155 2.13 ;
      RECT 0.96 0.625 1.69 0.955 ;
      RECT 1.485 2.13 1.655 2.3 ;
      RECT 1.405 2.3 1.655 2.735 ;
      RECT 0.115 2.475 0.365 2.98 ;
      RECT 0.115 2.305 1.235 2.475 ;
      RECT 1.065 2.475 1.235 2.905 ;
      RECT 1.065 2.905 2.185 3.075 ;
      RECT 1.855 2.3 2.185 2.905 ;
      RECT 3.425 2.12 3.675 2.98 ;
      RECT 3.425 1.95 4.235 2.12 ;
      RECT 4.065 1.67 4.235 1.95 ;
      RECT 4.065 1.34 4.445 1.67 ;
      RECT 4.065 1.17 4.235 1.34 ;
      RECT 3.42 1 4.235 1.17 ;
      RECT 2.945 1.81 3.195 2.98 ;
      RECT 2.605 1.48 3.195 1.81 ;
      RECT 2.94 0.595 3.195 1.48 ;
      RECT 5.385 2.905 7.825 3.075 ;
      RECT 6.9 2.9 7.825 2.905 ;
      RECT 5.385 2.18 5.555 2.905 ;
      RECT 6.9 2.73 8.045 2.9 ;
      RECT 5.035 2.01 5.555 2.18 ;
      RECT 7.875 2.295 8.045 2.73 ;
      RECT 5.035 1.83 5.365 2.01 ;
      RECT 7.875 2.125 9.235 2.295 ;
      RECT 8.905 2.295 9.235 2.98 ;
      RECT 8.905 2.12 9.235 2.125 ;
      RECT 7.875 1.115 8.045 2.125 ;
      RECT 8.905 1.95 9.945 2.12 ;
      RECT 7.875 0.945 8.28 1.115 ;
      RECT 9.615 1.58 9.945 1.95 ;
      RECT 7.95 0.605 8.28 0.945 ;
      RECT 10.305 2.27 10.635 2.98 ;
      RECT 10.305 2.1 10.91 2.27 ;
      RECT 10.74 1.92 10.91 2.1 ;
      RECT 10.74 1.75 11.75 1.92 ;
      RECT 11.58 1.92 12.665 2.09 ;
      RECT 11.555 1.11 11.725 1.75 ;
      RECT 12.495 1.89 12.665 1.92 ;
      RECT 10.94 0.94 11.725 1.11 ;
      RECT 12.495 1.72 13.365 1.89 ;
      RECT 10.94 0.85 11.11 0.94 ;
      RECT 13.035 1.47 13.365 1.72 ;
      RECT 9.96 0.6 11.11 0.85 ;
      RECT 13.185 2.505 14.655 2.675 ;
      RECT 14.485 1.76 14.655 2.505 ;
      RECT 14.485 1.43 14.815 1.76 ;
    LAYER mcon ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 12.155 1.58 12.325 1.75 ;
      RECT 10.235 1.21 10.405 1.38 ;
      RECT 9.275 1.58 9.445 1.75 ;
      RECT 5.915 1.21 6.085 1.38 ;
      RECT 17.915 -0.085 18.085 0.085 ;
      RECT 17.435 -0.085 17.605 0.085 ;
      RECT 16.955 -0.085 17.125 0.085 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 17.915 3.245 18.085 3.415 ;
      RECT 17.435 3.245 17.605 3.415 ;
      RECT 16.955 3.245 17.125 3.415 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.515 3.245 15.685 3.415 ;
    LAYER met1 ;
      RECT 5.855 1.365 6.145 1.41 ;
      RECT 5.855 1.225 10.465 1.365 ;
      RECT 10.175 1.365 10.465 1.41 ;
      RECT 5.855 1.18 6.145 1.225 ;
      RECT 10.175 1.18 10.465 1.225 ;
  END
END scs8ls_sdfbbn_2

MACRO scs8ls_sdfbbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 15.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.055 1.86 11.365 2.15 ;
        RECT 10.125 1.8 11.365 1.86 ;
        RECT 10.125 1.86 10.295 2.015 ;
        RECT 10.125 1.69 11.385 1.8 ;
        RECT 10.095 2.015 10.295 2.185 ;
        RECT 11.055 1.52 11.385 1.69 ;
        RECT 10.095 2.185 10.265 2.905 ;
        RECT 8.855 2.905 10.265 3.075 ;
        RECT 8.855 2.335 9.025 2.905 ;
        RECT 7.935 2.165 9.025 2.335 ;
        RECT 7.935 2.335 8.105 2.905 ;
        RECT 7.095 2.905 8.105 3.075 ;
        RECT 7.095 1.655 7.265 2.905 ;
        RECT 7.045 1.41 7.375 1.655 ;
    END
    ANTENNAGATEAREA 0.47 ;
  END SETB

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.43 1.18 3.76 1.67 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.395 0.35 15.735 2.98 ;
    END
    ANTENNADIFFAREA 0.5301 ;
  END Q

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.125 0.55 2.135 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805 1.55 1.285 2.095 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455 1.525 1.765 1.855 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.065 1.18 13.36 1.55 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END RESETB

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.87 1.72 14.275 2.89 ;
        RECT 14.105 1.05 14.275 1.72 ;
        RECT 13.77 0.35 14.275 1.05 ;
    END
    ANTENNADIFFAREA 0.5189 ;
  END QN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 15.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 15.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 12.635 1.21 12.805 1.38 ;
      RECT 8.315 1.21 8.485 1.38 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
    LAYER met1 ;
      RECT 8.255 1.365 8.545 1.41 ;
      RECT 8.255 1.225 12.865 1.365 ;
      RECT 12.575 1.365 12.865 1.41 ;
      RECT 8.255 1.18 8.545 1.225 ;
      RECT 12.575 1.18 12.865 1.225 ;
    LAYER li1 ;
      RECT 7.145 0.48 7.64 0.56 ;
      RECT 7.145 0.31 8.715 0.48 ;
      RECT 8.33 0.48 8.715 0.56 ;
      RECT 7.435 1.825 9.015 1.995 ;
      RECT 8.685 1.335 9.015 1.825 ;
      RECT 8.685 0.9 8.855 1.335 ;
      RECT 6.295 0.73 8.855 0.9 ;
      RECT 6.295 0.9 6.535 1.485 ;
      RECT 7.435 1.995 7.765 2.735 ;
      RECT 7.82 0.655 8.15 0.73 ;
      RECT 9.445 0.255 10.485 0.425 ;
      RECT 10.155 0.425 10.485 1.18 ;
      RECT 9.255 1.505 9.585 1.94 ;
      RECT 9.255 1.335 9.615 1.505 ;
      RECT 9.445 0.425 9.615 1.335 ;
      RECT 14.445 1.685 14.775 2.98 ;
      RECT 14.445 1.355 14.845 1.685 ;
      RECT 14.445 0.35 14.715 1.355 ;
      RECT 2.955 2.35 3.285 2.98 ;
      RECT 2.275 2.18 3.285 2.35 ;
      RECT 2.275 1.83 2.78 2.18 ;
      RECT 2.61 1.035 2.78 1.83 ;
      RECT 2.61 0.595 2.86 1.035 ;
      RECT 2.25 0.255 3.68 0.425 ;
      RECT 3.51 0.425 3.68 0.66 ;
      RECT 3.51 0.66 5.335 0.83 ;
      RECT 5.165 0.83 5.335 1.025 ;
      RECT 5.005 0.46 5.335 0.66 ;
      RECT 5.165 1.025 5.785 1.195 ;
      RECT 5.615 1.195 5.785 1.865 ;
      RECT 5.075 1.865 5.785 2.035 ;
      RECT 5.075 2.035 5.405 2.755 ;
      RECT 1.495 2.195 1.745 2.735 ;
      RECT 1.495 2.025 2.105 2.195 ;
      RECT 1.935 1.355 2.105 2.025 ;
      RECT 1.04 1.185 2.42 1.355 ;
      RECT 2.25 0.425 2.42 1.185 ;
      RECT 1.04 0.575 1.37 1.185 ;
      RECT 11.33 0.425 11.66 1.01 ;
      RECT 11.33 0.255 12.555 0.425 ;
      RECT 12.385 0.425 12.555 1.01 ;
      RECT 1.115 2.905 2.275 3.075 ;
      RECT 1.945 2.52 2.275 2.905 ;
      RECT 1.115 2.475 1.285 2.905 ;
      RECT 0.115 2.305 1.285 2.475 ;
      RECT 0.115 2.475 0.445 2.98 ;
      RECT 4.415 1.84 4.905 2.98 ;
      RECT 4.735 1.695 4.905 1.84 ;
      RECT 4.735 1.365 5.445 1.695 ;
      RECT 4.735 1.17 4.905 1.365 ;
      RECT 4.36 1 4.905 1.17 ;
      RECT 10.715 1.18 11.875 1.35 ;
      RECT 11.595 1.35 11.875 1.55 ;
      RECT 9.375 2.11 9.925 2.735 ;
      RECT 9.755 1.845 9.925 2.11 ;
      RECT 9.755 1.675 9.955 1.845 ;
      RECT 9.785 1.52 9.955 1.675 ;
      RECT 9.785 0.595 9.985 1.35 ;
      RECT 9.785 1.35 10.885 1.52 ;
      RECT 12.725 1.72 13.155 1.97 ;
      RECT 12.725 0.67 13.115 1.01 ;
      RECT 12.445 1.18 12.895 1.72 ;
      RECT 12.725 1.01 12.895 1.18 ;
      RECT 8.125 1.18 8.515 1.585 ;
      RECT 3.515 2.01 3.845 2.98 ;
      RECT 3.09 1.84 4.245 2.01 ;
      RECT 4.075 1.67 4.245 1.84 ;
      RECT 4.075 1.34 4.565 1.67 ;
      RECT 3.09 1.01 3.26 1.84 ;
      RECT 3.09 0.595 3.34 1.01 ;
      RECT 6.705 1.07 7.915 1.24 ;
      RECT 7.585 1.24 7.915 1.585 ;
      RECT 5.575 2.205 6.125 2.535 ;
      RECT 5.955 1.825 6.125 2.205 ;
      RECT 5.955 1.655 6.875 1.825 ;
      RECT 6.705 1.24 6.875 1.655 ;
      RECT 5.955 0.855 6.125 1.655 ;
      RECT 5.505 0.685 6.125 0.855 ;
      RECT 5.505 0.46 5.835 0.685 ;
      RECT 13.53 1.22 13.915 1.55 ;
      RECT 11.535 2.14 13.7 2.31 ;
      RECT 13.53 1.55 13.7 2.14 ;
      RECT 11.535 2.49 11.785 2.98 ;
      RECT 10.465 2.32 11.785 2.49 ;
      RECT 11.535 2.31 11.785 2.32 ;
      RECT 11.535 1.97 12.215 2.14 ;
      RECT 12.045 1.01 12.215 1.97 ;
      RECT 11.87 0.595 12.215 1.01 ;
      RECT 10.465 2.03 10.795 2.32 ;
      RECT 0 3.245 15.84 3.415 ;
      RECT 14.945 2.115 15.205 3.245 ;
      RECT 10.435 2.66 11.15 3.245 ;
      RECT 12.295 2.48 12.625 3.245 ;
      RECT 13.34 2.48 13.67 3.245 ;
      RECT 0.615 2.645 0.945 3.245 ;
      RECT 2.505 2.52 2.755 3.245 ;
      RECT 4.045 2.18 4.215 3.245 ;
      RECT 6.595 2.075 6.925 3.245 ;
      RECT 8.315 2.505 8.685 3.245 ;
      RECT 0 -0.085 15.84 0.085 ;
      RECT 14.895 0.085 15.225 0.94 ;
      RECT 0.14 0.085 0.47 0.955 ;
      RECT 1.83 0.085 2.08 1.015 ;
      RECT 3.85 0.085 4.18 0.49 ;
      RECT 6.49 0.085 6.885 0.56 ;
      RECT 9.025 0.085 9.275 1.05 ;
      RECT 10.9 0.085 11.15 1.01 ;
      RECT 13.295 0.085 13.59 1 ;
  END
END scs8ls_sdfbbp_1

MACRO scs8ls_sdfrbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 13.92 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.47 0.35 13.835 1.13 ;
        RECT 13.665 1.13 13.835 1.82 ;
        RECT 13.555 1.82 13.835 2.98 ;
    END
    ANTENNADIFFAREA 0.5189 LAYER met1 ;
    ANTENNADIFFAREA 0.5189 LAYER met2 ;
    ANTENNADIFFAREA 0.5189 LAYER met3 ;
    ANTENNADIFFAREA 0.5189 LAYER met4 ;
    ANTENNADIFFAREA 0.5189 LAYER met5 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.81 2.1 1.31 ;
    END
    ANTENNAGATEAREA 0.159 LAYER met1 ;
    ANTENNAGATEAREA 0.159 LAYER met2 ;
    ANTENNAGATEAREA 0.159 LAYER met3 ;
    ANTENNAGATEAREA 0.159 LAYER met4 ;
    ANTENNAGATEAREA 0.159 LAYER met5 ;
  END D

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.935 1.44 3.265 2.15 ;
    END
    ANTENNAGATEAREA 0.159 LAYER met1 ;
    ANTENNAGATEAREA 0.159 LAYER met2 ;
    ANTENNAGATEAREA 0.159 LAYER met3 ;
    ANTENNAGATEAREA 0.159 LAYER met4 ;
    ANTENNAGATEAREA 0.159 LAYER met5 ;
  END SCD

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.785 1.18 4.645 1.63 ;
        RECT 3.785 0.92 4.06 1.18 ;
    END
    ANTENNAGATEAREA 0.261 LAYER met1 ;
    ANTENNAGATEAREA 0.261 LAYER met2 ;
    ANTENNAGATEAREA 0.261 LAYER met3 ;
    ANTENNAGATEAREA 0.261 LAYER met4 ;
    ANTENNAGATEAREA 0.261 LAYER met5 ;
  END CLK

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.66 1.795 1.88 ;
        RECT 0.605 1.49 2.725 1.66 ;
        RECT 2.395 1.26 2.725 1.49 ;
    END
    ANTENNAGATEAREA 0.318 LAYER met1 ;
    ANTENNAGATEAREA 0.318 LAYER met2 ;
    ANTENNAGATEAREA 0.318 LAYER met3 ;
    ANTENNAGATEAREA 0.318 LAYER met4 ;
    ANTENNAGATEAREA 0.318 LAYER met5 ;
  END SCE

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.015 0.35 12.345 2.98 ;
    END
    ANTENNADIFFAREA 0.5376 LAYER met1 ;
    ANTENNADIFFAREA 0.5376 LAYER met2 ;
    ANTENNADIFFAREA 0.5376 LAYER met3 ;
    ANTENNADIFFAREA 0.5376 LAYER met4 ;
    ANTENNADIFFAREA 0.5376 LAYER met5 ;
  END QN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.92 3.575 ;
    END
  END vpwr

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3.935 1.965 10.945 2.105 ;
        RECT 10.655 2.105 10.945 2.15 ;
        RECT 10.655 1.92 10.945 1.965 ;
        RECT 3.935 2.105 4.225 2.15 ;
        RECT 7.775 2.105 8.065 2.15 ;
        RECT 3.935 1.92 4.225 1.965 ;
        RECT 7.775 1.92 8.065 1.965 ;
    END
    ANTENNAGATEAREA 0.411 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.956 LAYER met1 ;
    ANTENNAGATEAREA 0.411 LAYER met2 ;
    ANTENNAGATEAREA 0.411 LAYER met3 ;
    ANTENNAGATEAREA 0.411 LAYER met4 ;
    ANTENNAGATEAREA 0.411 LAYER met5 ;
  END RESETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 1.95 4.165 2.12 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 1.95 10.885 2.12 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 1.95 8.005 2.12 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
    LAYER li1 ;
      RECT 3.665 2.62 3.995 2.98 ;
      RECT 3.665 2.6 4.58 2.62 ;
      RECT 3.665 2.59 4.61 2.6 ;
      RECT 3.665 2.585 4.63 2.59 ;
      RECT 3.665 2.58 4.645 2.585 ;
      RECT 3.665 2.56 6.075 2.58 ;
      RECT 5.825 2.58 6.075 2.725 ;
      RECT 2.095 2.42 6.075 2.56 ;
      RECT 4.555 2.415 6.075 2.42 ;
      RECT 2.095 2.4 4.25 2.42 ;
      RECT 4.57 2.41 6.075 2.415 ;
      RECT 2.095 2.39 4.23 2.4 ;
      RECT 4.59 2.4 6.075 2.41 ;
      RECT 3.445 2.385 4.23 2.39 ;
      RECT 4.615 2.385 6.075 2.4 ;
      RECT 3.445 2.33 3.785 2.385 ;
      RECT 5.825 2.215 6.075 2.385 ;
      RECT 5.825 2.045 6.515 2.215 ;
      RECT 6.345 1.37 6.515 2.045 ;
      RECT 5.8 1.2 6.515 1.37 ;
      RECT 5.8 0.995 5.975 1.2 ;
      RECT 5.795 0.595 5.975 0.995 ;
      RECT 2.095 2.56 2.945 2.6 ;
      RECT 3.445 1.09 3.615 2.33 ;
      RECT 2.27 0.92 3.615 1.09 ;
      RECT 2.095 2.6 2.555 2.98 ;
      RECT 2.27 0.595 2.6 0.92 ;
      RECT 8.685 1.415 8.935 2.755 ;
      RECT 8.485 1.245 8.935 1.415 ;
      RECT 8.485 1.09 8.655 1.245 ;
      RECT 7.025 0.92 8.655 1.09 ;
      RECT 7.025 1.09 7.265 1.805 ;
      RECT 8.27 0.595 8.655 0.92 ;
      RECT 4.335 2.195 4.505 2.25 ;
      RECT 4.335 1.8 4.985 2.195 ;
      RECT 4.815 1.775 4.985 1.8 ;
      RECT 4.815 1.455 5.28 1.775 ;
      RECT 4.815 1.01 5.045 1.455 ;
      RECT 4.23 0.84 5.045 1.01 ;
      RECT 4.23 0.75 4.535 0.84 ;
      RECT 4.135 0.5 4.535 0.75 ;
      RECT 3.92 2.16 4.165 2.19 ;
      RECT 3.785 1.83 4.165 2.16 ;
      RECT 1.105 0.425 1.355 0.81 ;
      RECT 1.105 0.255 3.41 0.425 ;
      RECT 3.06 0.425 3.41 0.75 ;
      RECT 7.775 1.795 8.035 2.15 ;
      RECT 6.25 2.385 6.855 2.725 ;
      RECT 6.685 2.165 6.855 2.385 ;
      RECT 6.685 1.985 7.605 2.165 ;
      RECT 7.435 2.165 7.605 2.32 ;
      RECT 7.435 1.545 7.605 1.985 ;
      RECT 6.685 1.03 6.855 1.985 ;
      RECT 7.435 2.32 7.765 2.745 ;
      RECT 7.435 1.26 8.315 1.545 ;
      RECT 6.145 0.86 6.855 1.03 ;
      RECT 6.145 0.595 6.47 0.86 ;
      RECT 0 3.245 13.92 3.415 ;
      RECT 13.045 1.82 13.325 3.245 ;
      RECT 4.705 2.75 5.035 3.245 ;
      RECT 3.095 2.73 3.425 3.245 ;
      RECT 11.37 2.695 11.815 3.245 ;
      RECT 10.305 2.66 10.65 3.245 ;
      RECT 7.025 2.345 7.265 3.245 ;
      RECT 8.235 1.715 8.485 3.245 ;
      RECT 11.585 1.97 11.815 2.695 ;
      RECT 1.225 2.39 1.555 3.245 ;
      RECT 10.855 2.49 11.185 2.885 ;
      RECT 10.265 2.32 11.405 2.49 ;
      RECT 11.235 1.8 11.405 2.32 ;
      RECT 10.265 1.65 10.525 2.32 ;
      RECT 11.235 1.63 11.845 1.8 ;
      RECT 11.675 0.75 11.845 1.63 ;
      RECT 10.955 0.58 11.845 0.75 ;
      RECT 10.955 0.35 11.285 0.58 ;
      RECT 5.155 1.955 5.63 2.215 ;
      RECT 5.45 1.875 5.63 1.955 ;
      RECT 5.45 1.545 6.175 1.875 ;
      RECT 5.45 1.285 5.63 1.545 ;
      RECT 5.215 1.07 5.63 1.285 ;
      RECT 5.215 0.425 5.62 1.07 ;
      RECT 5.215 0.255 7.22 0.425 ;
      RECT 7.05 0.425 7.22 0.58 ;
      RECT 7.05 0.58 8.1 0.75 ;
      RECT 7.93 0.425 8.1 0.58 ;
      RECT 7.93 0.255 8.995 0.425 ;
      RECT 8.825 0.425 8.995 0.905 ;
      RECT 8.825 0.905 9.435 1.075 ;
      RECT 9.105 1.075 9.435 1.345 ;
      RECT 9.105 1.345 9.755 1.575 ;
      RECT 9.505 1.575 9.755 2.23 ;
      RECT 10.695 1.685 11.065 2.15 ;
      RECT 0.115 2.05 2.695 2.22 ;
      RECT 2.365 1.83 2.695 2.05 ;
      RECT 0.115 1.31 0.285 2.05 ;
      RECT 0.115 0.35 0.365 0.98 ;
      RECT 0.115 2.22 1.055 2.975 ;
      RECT 0.115 0.98 1.395 1.31 ;
      RECT 9.105 2.425 10.095 2.755 ;
      RECT 9.105 1.755 9.325 2.425 ;
      RECT 9.925 1.435 10.095 2.425 ;
      RECT 9.925 1.175 11.425 1.435 ;
      RECT 9.605 1.005 11.425 1.175 ;
      RECT 9.605 0.735 9.775 1.005 ;
      RECT 9.165 0.405 9.775 0.735 ;
      RECT 12.57 1.3 13.485 1.63 ;
      RECT 12.57 1.63 12.855 2.98 ;
      RECT 12.57 0.455 12.855 1.3 ;
      RECT 0 -0.085 13.92 0.085 ;
      RECT 13.12 0.085 13.29 1.13 ;
      RECT 3.59 0.085 3.88 0.75 ;
      RECT 4.705 0.085 5.035 0.67 ;
      RECT 7.43 0.085 7.76 0.41 ;
      RECT 10.165 0.085 10.495 0.76 ;
      RECT 11.51 0.085 11.84 0.41 ;
      RECT 0.545 0.085 0.875 0.81 ;
  END
END scs8ls_sdfrbp_1

MACRO scs8ls_sdfrbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 14.88 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.03 0.915 12.465 1.085 ;
        RECT 12.03 1.085 12.36 2.98 ;
        RECT 12.135 0.35 12.465 0.915 ;
    END
    ANTENNADIFFAREA 0.5432 LAYER met1 ;
    ANTENNADIFFAREA 0.5432 LAYER met2 ;
    ANTENNADIFFAREA 0.5432 LAYER met3 ;
    ANTENNADIFFAREA 0.5432 LAYER met4 ;
    ANTENNADIFFAREA 0.5432 LAYER met5 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.055 0.35 14.325 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 LAYER met1 ;
    ANTENNADIFFAREA 0.5432 LAYER met2 ;
    ANTENNADIFFAREA 0.5432 LAYER met3 ;
    ANTENNADIFFAREA 0.5432 LAYER met4 ;
    ANTENNADIFFAREA 0.5432 LAYER met5 ;
  END Q

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.945 1.44 3.275 2.15 ;
    END
    ANTENNAGATEAREA 0.159 LAYER met1 ;
    ANTENNAGATEAREA 0.159 LAYER met2 ;
    ANTENNAGATEAREA 0.159 LAYER met3 ;
    ANTENNAGATEAREA 0.159 LAYER met4 ;
    ANTENNAGATEAREA 0.159 LAYER met5 ;
  END SCD

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.54 1.82 1.795 2.15 ;
        RECT 1.625 1.62 1.795 1.82 ;
        RECT 1.625 1.36 2.735 1.62 ;
    END
    ANTENNAGATEAREA 0.318 LAYER met1 ;
    ANTENNAGATEAREA 0.318 LAYER met2 ;
    ANTENNAGATEAREA 0.318 LAYER met3 ;
    ANTENNAGATEAREA 0.318 LAYER met4 ;
    ANTENNAGATEAREA 0.318 LAYER met5 ;
  END SCE

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.905 1.18 4.235 1.55 ;
    END
    ANTENNAGATEAREA 0.261 LAYER met1 ;
    ANTENNAGATEAREA 0.261 LAYER met2 ;
    ANTENNAGATEAREA 0.261 LAYER met3 ;
    ANTENNAGATEAREA 0.261 LAYER met4 ;
    ANTENNAGATEAREA 0.261 LAYER met5 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.81 2.09 1.19 ;
    END
    ANTENNAGATEAREA 0.159 LAYER met1 ;
    ANTENNAGATEAREA 0.159 LAYER met2 ;
    ANTENNAGATEAREA 0.159 LAYER met3 ;
    ANTENNAGATEAREA 0.159 LAYER met4 ;
    ANTENNAGATEAREA 0.159 LAYER met5 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.88 3.575 ;
    END
  END vpwr

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3.935 1.965 10.945 2.105 ;
        RECT 3.935 2.105 4.225 2.15 ;
        RECT 7.775 2.105 8.065 2.15 ;
        RECT 10.655 2.105 10.945 2.15 ;
        RECT 3.935 1.92 4.225 1.965 ;
        RECT 7.775 1.92 8.065 1.965 ;
        RECT 10.655 1.92 10.945 1.965 ;
    END
    ANTENNAGATEAREA 0.411 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.956 LAYER met1 ;
    ANTENNAGATEAREA 0.411 LAYER met2 ;
    ANTENNAGATEAREA 0.411 LAYER met3 ;
    ANTENNAGATEAREA 0.411 LAYER met4 ;
    ANTENNAGATEAREA 0.411 LAYER met5 ;
  END RESETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 1.95 4.165 2.12 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 1.95 10.885 2.12 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 1.95 8.005 2.12 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
    LAYER li1 ;
      RECT 9.1 2.365 10.095 2.695 ;
      RECT 9.925 1.31 10.095 2.365 ;
      RECT 9.925 1.045 11.52 1.31 ;
      RECT 9.925 0.735 10.095 1.045 ;
      RECT 9.44 0.405 10.095 0.735 ;
      RECT 0 -0.085 14.88 0.085 ;
      RECT 14.495 0.085 14.78 1.13 ;
      RECT 12.635 0.085 12.895 1.05 ;
      RECT 13.67 0.085 13.84 1.13 ;
      RECT 3.64 0.085 3.97 0.835 ;
      RECT 4.75 0.085 4.92 1.13 ;
      RECT 7.45 0.085 7.985 0.41 ;
      RECT 10.335 0.085 10.665 0.81 ;
      RECT 11.645 0.085 11.895 0.535 ;
      RECT 0.545 0.085 0.875 0.835 ;
      RECT 10.715 1.82 11.395 2.15 ;
      RECT 5.155 2.03 5.63 2.24 ;
      RECT 5.155 1.985 5.675 2.03 ;
      RECT 5.155 1.945 6.15 1.985 ;
      RECT 5.43 1.9 6.15 1.945 ;
      RECT 5.475 1.5 6.15 1.9 ;
      RECT 5.475 1.275 5.645 1.5 ;
      RECT 5.1 0.99 5.645 1.275 ;
      RECT 5.1 0.48 5.43 0.99 ;
      RECT 5.1 0.31 7.17 0.48 ;
      RECT 7 0.48 7.17 0.58 ;
      RECT 7 0.58 8.325 0.75 ;
      RECT 8.155 0.425 8.325 0.58 ;
      RECT 8.155 0.255 9.27 0.425 ;
      RECT 9.1 0.425 9.27 0.905 ;
      RECT 9.1 0.905 9.64 1.235 ;
      RECT 9.31 1.235 9.64 1.865 ;
      RECT 9.31 1.865 9.755 2.195 ;
      RECT 8.64 1.745 8.93 2.755 ;
      RECT 8.76 1.09 8.93 1.745 ;
      RECT 7 0.92 8.93 1.09 ;
      RECT 7 1.09 7.21 1.78 ;
      RECT 8.495 0.595 8.93 0.92 ;
      RECT 6.16 2.51 6.9 2.725 ;
      RECT 6.16 2.495 7.915 2.51 ;
      RECT 7.55 2.51 7.915 2.725 ;
      RECT 6.66 2.34 7.915 2.495 ;
      RECT 7.38 2.32 7.915 2.34 ;
      RECT 6.66 0.95 6.83 2.34 ;
      RECT 7.38 1.575 7.55 2.32 ;
      RECT 6.16 0.65 6.83 0.95 ;
      RECT 7.38 1.26 8.59 1.575 ;
      RECT 7.72 1.795 8.02 2.15 ;
      RECT 2.775 2.42 5.985 2.49 ;
      RECT 3.615 2.49 5.985 2.58 ;
      RECT 4.57 2.41 5.985 2.42 ;
      RECT 2.775 2.32 3.995 2.42 ;
      RECT 3.615 2.58 4.645 2.59 ;
      RECT 5.71 2.58 5.985 2.725 ;
      RECT 5.8 2.325 5.985 2.41 ;
      RECT 3.615 2.59 3.995 2.98 ;
      RECT 5.8 2.155 6.49 2.325 ;
      RECT 6.32 1.29 6.49 2.155 ;
      RECT 5.82 1.12 6.49 1.29 ;
      RECT 5.82 0.82 5.99 1.12 ;
      RECT 5.66 0.65 5.99 0.82 ;
      RECT 1.94 2.66 2.945 2.91 ;
      RECT 2.775 2.49 2.945 2.66 ;
      RECT 3.445 1.175 3.615 2.32 ;
      RECT 2.26 1.005 3.615 1.175 ;
      RECT 2.26 0.595 2.61 1.005 ;
      RECT 13.065 1.63 13.325 2.98 ;
      RECT 13.065 1.3 13.885 1.63 ;
      RECT 13.065 0.35 13.325 1.3 ;
      RECT 4.335 1.99 4.505 2.25 ;
      RECT 4.335 1.82 4.985 1.99 ;
      RECT 4.405 1.775 4.985 1.82 ;
      RECT 4.405 1.445 5.305 1.775 ;
      RECT 4.405 1.01 4.575 1.445 ;
      RECT 4.24 0.595 4.575 1.01 ;
      RECT 11.065 2.49 11.395 2.795 ;
      RECT 10.265 2.32 11.395 2.49 ;
      RECT 10.265 1.65 10.545 2.32 ;
      RECT 10.265 1.48 11.86 1.65 ;
      RECT 11.69 0.875 11.86 1.48 ;
      RECT 11.125 0.705 11.86 0.875 ;
      RECT 11.125 0.35 11.455 0.705 ;
      RECT 0 3.245 14.88 3.415 ;
      RECT 14.495 1.82 14.775 3.245 ;
      RECT 12.54 1.92 12.83 3.245 ;
      RECT 13.545 1.82 13.875 3.245 ;
      RECT 4.705 2.75 5.035 3.245 ;
      RECT 7.07 2.68 7.32 3.245 ;
      RECT 3.115 2.66 3.445 3.245 ;
      RECT 10.265 2.66 10.86 3.245 ;
      RECT 11.6 1.82 11.85 3.245 ;
      RECT 8.19 1.745 8.44 3.245 ;
      RECT 0.615 2.73 1.4 3.245 ;
      RECT 3.785 1.82 4.165 2.15 ;
      RECT 1.095 0.255 3.43 0.425 ;
      RECT 3.1 0.425 3.43 0.835 ;
      RECT 1.095 0.425 1.345 0.835 ;
      RECT 0.115 2.32 2.605 2.49 ;
      RECT 2.275 1.83 2.605 2.32 ;
      RECT 0.115 2.49 0.445 2.98 ;
      RECT 0.115 1.58 0.285 2.32 ;
      RECT 0.115 0.375 0.365 1.25 ;
      RECT 0.115 1.25 1.395 1.58 ;
  END
END scs8ls_sdfrbp_2

MACRO scs8ls_sdfrtn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 13.92 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.78 1.98 2.12 ;
    END
    ANTENNAGATEAREA 0.159 LAYER met1 ;
    ANTENNAGATEAREA 0.159 LAYER met2 ;
    ANTENNAGATEAREA 0.159 LAYER met3 ;
    ANTENNAGATEAREA 0.159 LAYER met4 ;
    ANTENNAGATEAREA 0.159 LAYER met5 ;
  END D

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.875 0.955 2.55 1.41 ;
        RECT 0.535 1.41 2.045 1.58 ;
        RECT 0.535 1.58 0.865 2.08 ;
    END
    ANTENNAGATEAREA 0.318 LAYER met1 ;
    ANTENNAGATEAREA 0.318 LAYER met2 ;
    ANTENNAGATEAREA 0.318 LAYER met3 ;
    ANTENNAGATEAREA 0.318 LAYER met4 ;
    ANTENNAGATEAREA 0.318 LAYER met5 ;
  END SCE

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.8 1.525 3.235 2.15 ;
    END
    ANTENNAGATEAREA 0.159 LAYER met1 ;
    ANTENNAGATEAREA 0.159 LAYER met2 ;
    ANTENNAGATEAREA 0.159 LAYER met3 ;
    ANTENNAGATEAREA 0.159 LAYER met4 ;
    ANTENNAGATEAREA 0.159 LAYER met5 ;
  END SCD

  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.275 1.21 4.675 1.55 ;
    END
    ANTENNAGATEAREA 0.261 LAYER met1 ;
    ANTENNAGATEAREA 0.261 LAYER met2 ;
    ANTENNAGATEAREA 0.261 LAYER met3 ;
    ANTENNAGATEAREA 0.261 LAYER met4 ;
    ANTENNAGATEAREA 0.261 LAYER met5 ;
  END CLKN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.475 0.35 13.805 2.98 ;
    END
    ANTENNADIFFAREA 0.5469 LAYER met1 ;
    ANTENNADIFFAREA 0.5469 LAYER met2 ;
    ANTENNADIFFAREA 0.5469 LAYER met3 ;
    ANTENNADIFFAREA 0.5469 LAYER met4 ;
    ANTENNADIFFAREA 0.5469 LAYER met5 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.92 3.575 ;
    END
  END vpwr

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3.455 1.595 11.425 1.735 ;
        RECT 3.455 1.735 3.745 1.78 ;
        RECT 3.455 1.55 3.745 1.595 ;
        RECT 7.775 1.735 8.065 1.78 ;
        RECT 11.135 1.735 11.425 1.78 ;
        RECT 7.775 1.55 8.065 1.595 ;
        RECT 11.135 1.55 11.425 1.595 ;
    END
    ANTENNAGATEAREA 0.411 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 5.628 LAYER met1 ;
    ANTENNAGATEAREA 0.411 LAYER met2 ;
    ANTENNAGATEAREA 0.411 LAYER met3 ;
    ANTENNAGATEAREA 0.411 LAYER met4 ;
    ANTENNAGATEAREA 0.411 LAYER met5 ;
  END RESETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 1.58 8.005 1.75 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 1.58 3.685 1.75 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 1.58 11.365 1.75 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
    LAYER li1 ;
      RECT 9.03 1.54 9.35 1.8 ;
      RECT 9.03 1.47 10.395 1.54 ;
      RECT 9.18 1.37 10.395 1.47 ;
      RECT 10.065 1.225 10.395 1.37 ;
      RECT 6.495 1.99 6.715 2.065 ;
      RECT 5.23 1.775 6.715 1.99 ;
      RECT 5.425 1.735 6.715 1.775 ;
      RECT 5.425 1.465 5.675 1.735 ;
      RECT 5.425 1.265 6.495 1.465 ;
      RECT 5.425 1.085 5.675 1.265 ;
      RECT 6.325 0.545 6.495 1.265 ;
      RECT 5.345 0.87 5.675 1.085 ;
      RECT 6.325 0.255 7.72 0.545 ;
      RECT 7.495 0.545 7.72 0.79 ;
      RECT 7.495 0.79 9.825 0.96 ;
      RECT 9.495 0.96 9.825 1.2 ;
      RECT 8.795 2.14 9.565 2.98 ;
      RECT 8.69 1.97 9.565 2.14 ;
      RECT 8.69 1.3 8.86 1.97 ;
      RECT 7.225 1.13 9.01 1.3 ;
      RECT 7.225 1.3 7.475 1.87 ;
      RECT 6.285 2.445 6.57 2.735 ;
      RECT 6.285 2.235 7.055 2.445 ;
      RECT 6.885 2.21 7.055 2.235 ;
      RECT 6.885 2.14 7.95 2.21 ;
      RECT 7.575 2.21 7.95 2.735 ;
      RECT 6.885 2.04 8.52 2.14 ;
      RECT 7.645 1.97 8.52 2.04 ;
      RECT 6.885 1.095 7.055 2.04 ;
      RECT 8.225 1.47 8.52 1.97 ;
      RECT 6.665 0.725 7.055 1.095 ;
      RECT 7.685 1.47 8.035 1.8 ;
      RECT 3.43 2.35 4.645 2.395 ;
      RECT 3.43 2.34 4.7 2.35 ;
      RECT 3.43 2.33 4.72 2.34 ;
      RECT 3.43 2.195 6.115 2.33 ;
      RECT 5.855 2.33 6.115 2.735 ;
      RECT 3.905 2.17 6.115 2.195 ;
      RECT 4.66 2.16 6.115 2.17 ;
      RECT 3.905 0.53 6.155 0.7 ;
      RECT 5.905 0.7 6.155 1.095 ;
      RECT 1.405 2.63 3.68 2.8 ;
      RECT 3.43 2.8 3.68 2.98 ;
      RECT 3.43 2.395 3.68 2.63 ;
      RECT 3.905 1.185 4.075 2.17 ;
      RECT 2.72 1.015 4.075 1.185 ;
      RECT 2.72 0.765 2.89 1.015 ;
      RECT 3.905 0.7 4.075 1.015 ;
      RECT 1.955 0.595 2.89 0.765 ;
      RECT 1.405 2.8 2.22 2.96 ;
      RECT 4.255 1.99 4.6 2 ;
      RECT 4.255 1.82 5.03 1.99 ;
      RECT 4.845 1.605 5.03 1.82 ;
      RECT 4.845 1.235 5.255 1.605 ;
      RECT 4.845 1.04 5.165 1.235 ;
      RECT 4.245 0.87 5.165 1.04 ;
      RECT 0 3.245 13.92 3.415 ;
      RECT 2.815 2.97 3.145 3.245 ;
      RECT 10.605 2.65 11.21 3.245 ;
      RECT 11.88 2.63 12.21 3.245 ;
      RECT 4.78 2.5 5.11 3.245 ;
      RECT 7.225 2.38 7.395 3.245 ;
      RECT 8.295 2.31 8.625 3.245 ;
      RECT 12.975 1.82 13.305 3.245 ;
      RECT 0.565 2.63 0.895 3.245 ;
      RECT 11.195 1.54 11.395 1.78 ;
      RECT 10.995 1.21 11.395 1.54 ;
      RECT 9.735 1.88 10.065 2.98 ;
      RECT 9.735 1.71 11.025 1.88 ;
      RECT 10.855 1.88 11.025 1.95 ;
      RECT 10.855 1.95 11.895 2.12 ;
      RECT 11.565 1.04 11.895 1.95 ;
      RECT 9.995 0.87 11.895 1.04 ;
      RECT 9.995 0.62 10.165 0.87 ;
      RECT 9.19 0.29 10.165 0.62 ;
      RECT 11.38 2.46 11.71 2.98 ;
      RECT 10.435 2.29 12.235 2.46 ;
      RECT 10.435 2.05 10.685 2.29 ;
      RECT 12.065 0.7 12.235 2.29 ;
      RECT 11.69 0.45 12.235 0.7 ;
      RECT 12.44 1.685 12.795 2.98 ;
      RECT 12.44 1.355 12.81 1.685 ;
      RECT 12.44 0.35 12.795 1.355 ;
      RECT 0 -0.085 13.92 0.085 ;
      RECT 3.575 0.085 4.065 0.36 ;
      RECT 4.805 0.085 5.165 0.36 ;
      RECT 7.89 0.085 8.22 0.62 ;
      RECT 10.73 0.085 11.2 0.68 ;
      RECT 12.975 0.085 13.305 1.13 ;
      RECT 0.615 0.085 0.945 0.88 ;
      RECT 3.405 1.355 3.735 2.025 ;
      RECT 1.165 0.425 1.495 0.765 ;
      RECT 1.165 0.255 3.39 0.425 ;
      RECT 3.06 0.425 3.39 0.845 ;
      RECT 0.115 2.29 2.545 2.46 ;
      RECT 2.215 1.58 2.545 2.29 ;
      RECT 0.115 2.46 0.365 2.98 ;
      RECT 0.115 1.24 0.365 2.29 ;
      RECT 0.115 0.42 0.445 1.05 ;
      RECT 0.115 1.05 1.62 1.24 ;
      RECT 1.29 0.935 1.62 1.05 ;
  END
END scs8ls_sdfrtn_1

MACRO scs8ls_sdfrtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.81 2.1 1.265 ;
    END
    ANTENNAGATEAREA 0.159 LAYER met1 ;
    ANTENNAGATEAREA 0.159 LAYER met2 ;
    ANTENNAGATEAREA 0.159 LAYER met3 ;
    ANTENNAGATEAREA 0.159 LAYER met4 ;
    ANTENNAGATEAREA 0.159 LAYER met5 ;
  END D

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.945 1.44 3.275 2.15 ;
    END
    ANTENNAGATEAREA 0.159 LAYER met1 ;
    ANTENNAGATEAREA 0.159 LAYER met2 ;
    ANTENNAGATEAREA 0.159 LAYER met3 ;
    ANTENNAGATEAREA 0.159 LAYER met4 ;
    ANTENNAGATEAREA 0.159 LAYER met5 ;
  END SCD

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.785 1.26 4.64 1.65 ;
        RECT 3.785 0.92 4.195 1.26 ;
    END
    ANTENNAGATEAREA 0.261 LAYER met1 ;
    ANTENNAGATEAREA 0.261 LAYER met2 ;
    ANTENNAGATEAREA 0.261 LAYER met3 ;
    ANTENNAGATEAREA 0.261 LAYER met4 ;
    ANTENNAGATEAREA 0.261 LAYER met5 ;
  END CLK

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455 1.66 1.795 1.835 ;
        RECT 0.455 1.49 2.725 1.66 ;
        RECT 2.345 1.26 2.725 1.49 ;
    END
    ANTENNAGATEAREA 0.318 LAYER met1 ;
    ANTENNAGATEAREA 0.318 LAYER met2 ;
    ANTENNAGATEAREA 0.318 LAYER met3 ;
    ANTENNAGATEAREA 0.318 LAYER met4 ;
    ANTENNAGATEAREA 0.318 LAYER met5 ;
  END SCE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.995 0.35 13.325 1.13 ;
        RECT 13.07 1.13 13.325 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 LAYER met1 ;
    ANTENNADIFFAREA 0.5413 LAYER met2 ;
    ANTENNADIFFAREA 0.5413 LAYER met3 ;
    ANTENNADIFFAREA 0.5413 LAYER met4 ;
    ANTENNADIFFAREA 0.5413 LAYER met5 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.44 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.44 3.575 ;
    END
  END vpwr

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3.935 1.965 10.945 2.105 ;
        RECT 10.655 2.105 10.945 2.15 ;
        RECT 10.655 1.92 10.945 1.965 ;
        RECT 3.935 2.105 4.225 2.15 ;
        RECT 7.775 2.105 8.065 2.15 ;
        RECT 3.935 1.92 4.225 1.965 ;
        RECT 7.775 1.92 8.065 1.965 ;
    END
    ANTENNAGATEAREA 0.411 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.956 LAYER met1 ;
    ANTENNAGATEAREA 0.411 LAYER met2 ;
    ANTENNAGATEAREA 0.411 LAYER met3 ;
    ANTENNAGATEAREA 0.411 LAYER met4 ;
    ANTENNAGATEAREA 0.411 LAYER met5 ;
  END RESETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 1.95 8.005 2.12 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 1.95 4.165 2.12 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 1.95 10.885 2.12 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
    LAYER li1 ;
      RECT 0 -0.085 13.44 0.085 ;
      RECT 3.59 0.085 3.88 0.75 ;
      RECT 4.705 0.085 5.035 0.75 ;
      RECT 7.43 0.085 7.76 0.41 ;
      RECT 10.195 0.085 10.525 0.81 ;
      RECT 11.57 0.085 11.905 0.585 ;
      RECT 12.565 0.085 12.815 1.13 ;
      RECT 0.545 0.085 0.875 0.88 ;
      RECT 0 3.245 13.44 3.415 ;
      RECT 4.705 2.75 5.035 3.245 ;
      RECT 3.095 2.685 3.425 3.245 ;
      RECT 7.205 2.66 7.54 3.245 ;
      RECT 10.485 2.52 10.735 3.245 ;
      RECT 11.48 2.1 11.81 3.245 ;
      RECT 12.54 1.82 12.87 3.245 ;
      RECT 8.385 1.745 8.555 3.245 ;
      RECT 0.615 2.345 0.945 3.245 ;
      RECT 11.98 2.1 12.31 2.98 ;
      RECT 12.085 1.63 12.31 2.1 ;
      RECT 12.085 1.3 12.87 1.63 ;
      RECT 12.085 0.35 12.335 1.3 ;
      RECT 10.945 2.52 11.31 2.98 ;
      RECT 11.14 1.615 11.31 2.52 ;
      RECT 9.985 1.445 11.735 1.615 ;
      RECT 9.985 1.435 10.315 1.445 ;
      RECT 11.565 0.925 11.735 1.445 ;
      RECT 11.01 0.755 11.735 0.925 ;
      RECT 11.01 0.35 11.34 0.755 ;
      RECT 9.29 2.55 10.315 2.88 ;
      RECT 10.145 1.955 10.315 2.55 ;
      RECT 9.585 1.785 10.315 1.955 ;
      RECT 9.585 1.265 9.755 1.785 ;
      RECT 9.585 1.095 11.395 1.265 ;
      RECT 11.065 1.265 11.395 1.275 ;
      RECT 9.585 0.77 9.755 1.095 ;
      RECT 9.405 0.35 9.755 0.77 ;
      RECT 10.64 1.82 10.97 2.15 ;
      RECT 9.245 2.125 9.975 2.38 ;
      RECT 9.245 1.27 9.415 2.125 ;
      RECT 9.065 0.94 9.415 1.27 ;
      RECT 9.065 0.425 9.235 0.94 ;
      RECT 7.93 0.255 9.235 0.425 ;
      RECT 7.93 0.425 8.1 0.58 ;
      RECT 7.05 0.58 8.1 0.75 ;
      RECT 7.05 0.425 7.22 0.58 ;
      RECT 5.215 0.255 7.22 0.425 ;
      RECT 5.215 0.425 5.62 1.07 ;
      RECT 5.215 1.07 5.63 1.285 ;
      RECT 5.45 1.285 5.63 1.545 ;
      RECT 5.45 1.545 6.2 1.875 ;
      RECT 5.45 1.875 5.63 1.955 ;
      RECT 5.155 1.955 5.63 2.215 ;
      RECT 8.725 1.715 9.005 2.755 ;
      RECT 8.725 1.09 8.895 1.715 ;
      RECT 7.05 0.92 8.895 1.09 ;
      RECT 7.05 1.09 7.325 1.805 ;
      RECT 8.27 0.595 8.655 0.92 ;
      RECT 6.25 2.49 6.88 2.725 ;
      RECT 6.25 2.385 8.075 2.49 ;
      RECT 7.745 2.49 8.075 2.745 ;
      RECT 6.71 2.32 8.075 2.385 ;
      RECT 7.495 1.575 7.665 2.32 ;
      RECT 6.71 1.03 6.88 2.32 ;
      RECT 7.495 1.26 8.315 1.575 ;
      RECT 6.145 0.86 6.88 1.03 ;
      RECT 6.145 0.595 6.47 0.86 ;
      RECT 7.835 1.815 8.165 2.15 ;
      RECT 3.665 2.62 3.995 2.98 ;
      RECT 3.665 2.6 4.58 2.62 ;
      RECT 3.665 2.59 4.61 2.6 ;
      RECT 3.665 2.585 4.63 2.59 ;
      RECT 3.665 2.58 4.645 2.585 ;
      RECT 3.665 2.515 6.075 2.58 ;
      RECT 5.825 2.58 6.075 2.725 ;
      RECT 1.485 2.42 6.075 2.515 ;
      RECT 4.555 2.415 6.075 2.42 ;
      RECT 1.485 2.4 4.25 2.42 ;
      RECT 4.57 2.41 6.075 2.415 ;
      RECT 1.485 2.385 4.23 2.4 ;
      RECT 4.59 2.4 6.075 2.41 ;
      RECT 1.485 2.345 3.785 2.385 ;
      RECT 4.615 2.385 6.075 2.4 ;
      RECT 3.445 2.33 3.785 2.345 ;
      RECT 5.825 2.215 6.075 2.385 ;
      RECT 5.825 2.045 6.54 2.215 ;
      RECT 6.37 1.37 6.54 2.045 ;
      RECT 5.8 1.2 6.54 1.37 ;
      RECT 5.8 0.995 5.975 1.2 ;
      RECT 5.795 0.595 5.975 0.995 ;
      RECT 3.445 1.09 3.615 2.33 ;
      RECT 2.27 0.92 3.615 1.09 ;
      RECT 1.485 2.515 2.555 2.98 ;
      RECT 2.27 0.595 2.6 0.92 ;
      RECT 4.335 2.195 4.505 2.25 ;
      RECT 4.335 1.82 4.98 2.195 ;
      RECT 4.81 1.775 4.98 1.82 ;
      RECT 4.81 1.455 5.28 1.775 ;
      RECT 4.81 1.09 5.045 1.455 ;
      RECT 4.365 0.92 5.045 1.09 ;
      RECT 4.365 0.75 4.535 0.92 ;
      RECT 4.135 0.5 4.535 0.75 ;
      RECT 3.92 2.16 4.165 2.19 ;
      RECT 3.785 1.83 4.165 2.16 ;
      RECT 1.105 0.425 1.435 0.64 ;
      RECT 1.105 0.255 3.41 0.425 ;
      RECT 3.06 0.425 3.41 0.75 ;
      RECT 0.115 2.005 2.705 2.175 ;
      RECT 2.035 1.83 2.705 2.005 ;
      RECT 0.115 2.175 0.445 2.98 ;
      RECT 0.115 1.265 0.285 2.005 ;
      RECT 0.115 0.42 0.365 1.05 ;
      RECT 0.115 1.05 1.375 1.265 ;
      RECT 1.045 0.935 1.375 1.05 ;
  END
END scs8ls_sdfrtp_1

MACRO scs8ls_sdfrtp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 14.4 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.525 0.35 13.855 1.41 ;
        RECT 13.525 1.41 13.785 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 LAYER met1 ;
    ANTENNADIFFAREA 0.5432 LAYER met2 ;
    ANTENNADIFFAREA 0.5432 LAYER met3 ;
    ANTENNADIFFAREA 0.5432 LAYER met4 ;
    ANTENNADIFFAREA 0.5432 LAYER met5 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.785 1.26 4.645 1.63 ;
        RECT 3.785 1.18 4.195 1.26 ;
        RECT 3.785 0.92 4.06 1.18 ;
    END
    ANTENNAGATEAREA 0.261 LAYER met1 ;
    ANTENNAGATEAREA 0.261 LAYER met2 ;
    ANTENNAGATEAREA 0.261 LAYER met3 ;
    ANTENNAGATEAREA 0.261 LAYER met4 ;
    ANTENNAGATEAREA 0.261 LAYER met5 ;
  END CLK

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.945 1.44 3.275 2 ;
        RECT 2.875 2 3.275 2.175 ;
    END
    ANTENNAGATEAREA 0.159 LAYER met1 ;
    ANTENNAGATEAREA 0.159 LAYER met2 ;
    ANTENNAGATEAREA 0.159 LAYER met3 ;
    ANTENNAGATEAREA 0.159 LAYER met4 ;
    ANTENNAGATEAREA 0.159 LAYER met5 ;
  END SCD

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455 1.66 2.205 1.835 ;
        RECT 0.455 1.49 2.705 1.66 ;
        RECT 2.375 1.26 2.705 1.49 ;
    END
    ANTENNAGATEAREA 0.318 LAYER met1 ;
    ANTENNAGATEAREA 0.318 LAYER met2 ;
    ANTENNAGATEAREA 0.318 LAYER met3 ;
    ANTENNAGATEAREA 0.318 LAYER met4 ;
    ANTENNAGATEAREA 0.318 LAYER met5 ;
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.81 2.1 1.265 ;
        RECT 1.605 0.595 2.1 0.81 ;
    END
    ANTENNAGATEAREA 0.159 LAYER met1 ;
    ANTENNAGATEAREA 0.159 LAYER met2 ;
    ANTENNAGATEAREA 0.159 LAYER met3 ;
    ANTENNAGATEAREA 0.159 LAYER met4 ;
    ANTENNAGATEAREA 0.159 LAYER met5 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.4 3.575 ;
    END
  END vpwr

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3.935 1.965 11.425 2.105 ;
        RECT 11.135 2.105 11.425 2.15 ;
        RECT 11.135 1.92 11.425 1.965 ;
        RECT 3.935 2.105 4.225 2.15 ;
        RECT 8.255 2.105 8.545 2.15 ;
        RECT 3.935 1.92 4.225 1.965 ;
        RECT 8.255 1.92 8.545 1.965 ;
    END
    ANTENNAGATEAREA 0.411 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 5.292 LAYER met1 ;
    ANTENNAGATEAREA 0.411 LAYER met2 ;
    ANTENNAGATEAREA 0.411 LAYER met3 ;
    ANTENNAGATEAREA 0.411 LAYER met4 ;
    ANTENNAGATEAREA 0.411 LAYER met5 ;
  END RESETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 7.435 1.545 7.605 1.985 ;
      RECT 6.685 1.03 6.855 1.985 ;
      RECT 7.435 2.32 7.765 2.745 ;
      RECT 7.435 1.26 8.485 1.545 ;
      RECT 6.145 0.86 6.855 1.03 ;
      RECT 6.145 0.595 6.47 0.86 ;
      RECT 11.41 2.56 11.74 2.98 ;
      RECT 10.56 2.39 11.74 2.56 ;
      RECT 10.56 1.75 10.85 2.39 ;
      RECT 10.56 1.58 12.23 1.75 ;
      RECT 10.56 1.37 10.85 1.58 ;
      RECT 12.06 0.94 12.23 1.58 ;
      RECT 11.545 0.77 12.23 0.94 ;
      RECT 11.545 0.35 11.875 0.77 ;
      RECT 0 3.245 14.4 3.415 ;
      RECT 13.955 1.82 14.285 3.245 ;
      RECT 4.705 2.75 5.035 3.245 ;
      RECT 10.56 2.73 11.24 3.245 ;
      RECT 3.095 2.685 3.425 3.245 ;
      RECT 7.025 2.345 7.265 3.245 ;
      RECT 8.245 2.33 8.58 3.245 ;
      RECT 11.945 1.94 12.275 3.245 ;
      RECT 13.005 1.82 13.335 3.245 ;
      RECT 0.615 2.345 1.565 3.245 ;
      RECT 12.445 1.94 12.775 2.98 ;
      RECT 12.605 1.63 12.775 1.94 ;
      RECT 12.605 1.3 13.355 1.63 ;
      RECT 12.605 0.35 12.865 1.3 ;
      RECT 11.11 1.92 11.44 2.22 ;
      RECT 8.75 1.715 9.115 2.755 ;
      RECT 8.75 1.09 8.92 1.715 ;
      RECT 7.025 0.92 8.92 1.09 ;
      RECT 7.025 1.09 7.265 1.805 ;
      RECT 8.27 0.595 8.92 0.92 ;
      RECT 7.775 1.795 8.57 2.15 ;
      RECT 4.335 2.195 4.505 2.25 ;
      RECT 4.335 1.82 4.985 2.195 ;
      RECT 4.815 1.775 4.985 1.82 ;
      RECT 4.815 1.455 5.28 1.775 ;
      RECT 4.815 1.08 5.045 1.455 ;
      RECT 4.39 0.935 5.045 1.08 ;
      RECT 4.37 0.91 5.045 0.935 ;
      RECT 4.355 0.89 5.045 0.91 ;
      RECT 4.345 0.88 5.045 0.89 ;
      RECT 4.325 0.865 4.625 0.88 ;
      RECT 4.3 0.86 4.625 0.865 ;
      RECT 4.3 0.845 4.6 0.86 ;
      RECT 4.23 0.835 4.58 0.845 ;
      RECT 4.23 0.815 4.57 0.835 ;
      RECT 4.23 0.79 4.555 0.815 ;
      RECT 4.23 0.75 4.535 0.79 ;
      RECT 4.135 0.5 4.535 0.75 ;
      RECT 0 -0.085 14.4 0.085 ;
      RECT 14.035 0.085 14.285 1.13 ;
      RECT 3.61 0.085 3.88 0.73 ;
      RECT 4.705 0.085 5.035 0.71 ;
      RECT 7.43 0.085 7.76 0.41 ;
      RECT 10.755 0.085 11.085 0.81 ;
      RECT 12.105 0.085 12.435 0.6 ;
      RECT 13.095 0.085 13.345 1.13 ;
      RECT 0.545 0.085 0.875 0.765 ;
      RECT 3.615 2.62 3.995 2.98 ;
      RECT 3.615 2.6 4.58 2.62 ;
      RECT 3.615 2.59 4.61 2.6 ;
      RECT 3.615 2.585 4.63 2.59 ;
      RECT 3.615 2.58 4.645 2.585 ;
      RECT 3.615 2.515 6.075 2.58 ;
      RECT 5.825 2.58 6.075 2.725 ;
      RECT 2.095 2.42 6.075 2.515 ;
      RECT 4.555 2.415 6.075 2.42 ;
      RECT 2.095 2.4 4.25 2.42 ;
      RECT 4.57 2.41 6.075 2.415 ;
      RECT 2.095 2.385 4.23 2.4 ;
      RECT 4.59 2.4 6.075 2.41 ;
      RECT 2.095 2.345 3.785 2.385 ;
      RECT 4.615 2.385 6.075 2.4 ;
      RECT 3.445 2.33 3.785 2.345 ;
      RECT 5.825 2.215 6.075 2.385 ;
      RECT 5.825 2.045 6.515 2.215 ;
      RECT 6.345 1.37 6.515 2.045 ;
      RECT 5.8 1.2 6.515 1.37 ;
      RECT 5.8 0.995 5.975 1.2 ;
      RECT 5.795 0.595 5.975 0.995 ;
      RECT 3.445 1.27 3.615 2.33 ;
      RECT 2.875 0.935 3.615 1.27 ;
      RECT 2.855 0.91 3.615 0.935 ;
      RECT 2.84 0.9 3.615 0.91 ;
      RECT 2.84 0.89 3.11 0.9 ;
      RECT 2.83 0.88 3.11 0.89 ;
      RECT 2.81 0.865 3.085 0.88 ;
      RECT 2.785 0.855 3.065 0.865 ;
      RECT 2.785 0.845 3.055 0.855 ;
      RECT 2.27 0.835 3.055 0.845 ;
      RECT 2.27 0.81 3.04 0.835 ;
      RECT 2.27 0.595 3.02 0.81 ;
      RECT 2.095 2.515 2.425 2.98 ;
      RECT 0.115 2.005 2.705 2.175 ;
      RECT 2.375 1.83 2.705 2.005 ;
      RECT 0.115 2.175 0.445 2.98 ;
      RECT 0.115 1.265 0.285 2.005 ;
      RECT 0.115 0.35 0.365 0.935 ;
      RECT 0.115 0.935 1.14 1.265 ;
      RECT 9.32 2.52 10.39 2.85 ;
      RECT 9.32 1.84 9.6 2.52 ;
      RECT 10.22 1.2 10.39 2.52 ;
      RECT 10.22 1.11 11.89 1.2 ;
      RECT 11.02 1.2 11.89 1.41 ;
      RECT 10.22 1.03 11.19 1.11 ;
      RECT 10.22 0.81 10.39 1.03 ;
      RECT 9.43 0.48 10.39 0.81 ;
      RECT 3.92 2.16 4.165 2.19 ;
      RECT 3.785 1.83 4.165 2.16 ;
      RECT 1.105 0.255 3.43 0.425 ;
      RECT 3.19 0.425 3.43 0.73 ;
      RECT 1.105 0.425 1.435 0.64 ;
      RECT 5.155 1.955 5.63 2.215 ;
      RECT 5.45 1.875 5.63 1.955 ;
      RECT 5.45 1.545 6.175 1.875 ;
      RECT 5.45 1.285 5.63 1.545 ;
      RECT 5.215 1.07 5.63 1.285 ;
      RECT 5.215 0.425 5.62 1.07 ;
      RECT 5.215 0.255 7.22 0.425 ;
      RECT 7.05 0.425 7.22 0.58 ;
      RECT 7.05 0.58 8.1 0.75 ;
      RECT 7.93 0.425 8.1 0.58 ;
      RECT 7.93 0.255 9.26 0.425 ;
      RECT 9.09 0.425 9.26 1.005 ;
      RECT 9.09 1.005 10.05 1.335 ;
      RECT 9.785 1.335 10.05 2.33 ;
      RECT 6.25 2.385 6.855 2.725 ;
      RECT 6.685 2.165 6.855 2.385 ;
      RECT 6.685 1.985 7.605 2.165 ;
      RECT 7.435 2.165 7.605 2.32 ;
    LAYER mcon ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 1.95 11.365 2.12 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 1.95 8.485 2.12 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 1.95 4.165 2.12 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_sdfrtp_2

MACRO scs8ls_sdfrtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 14.88 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.085 1.3 14.755 1.77 ;
        RECT 13.085 1.77 14.755 1.94 ;
        RECT 14.085 1.1 14.255 1.3 ;
        RECT 13.085 1.94 13.415 2.98 ;
        RECT 14.065 1.94 14.28 2.98 ;
        RECT 12.535 0.93 14.255 1.1 ;
        RECT 12.535 0.35 12.865 0.93 ;
        RECT 14.085 0.35 14.255 0.93 ;
    END
    ANTENNADIFFAREA 1.0864 LAYER met1 ;
    ANTENNADIFFAREA 1.0864 LAYER met2 ;
    ANTENNADIFFAREA 1.0864 LAYER met3 ;
    ANTENNADIFFAREA 1.0864 LAYER met4 ;
    ANTENNADIFFAREA 1.0864 LAYER met5 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.84 1.26 4.635 1.59 ;
        RECT 3.84 1.18 4.195 1.26 ;
    END
    ANTENNAGATEAREA 0.261 LAYER met1 ;
    ANTENNAGATEAREA 0.261 LAYER met2 ;
    ANTENNAGATEAREA 0.261 LAYER met3 ;
    ANTENNAGATEAREA 0.261 LAYER met4 ;
    ANTENNAGATEAREA 0.261 LAYER met5 ;
  END CLK

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.945 1.44 3.275 2.15 ;
    END
    ANTENNAGATEAREA 0.159 LAYER met1 ;
    ANTENNAGATEAREA 0.159 LAYER met2 ;
    ANTENNAGATEAREA 0.159 LAYER met3 ;
    ANTENNAGATEAREA 0.159 LAYER met4 ;
    ANTENNAGATEAREA 0.159 LAYER met5 ;
  END SCD

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.66 1.795 1.835 ;
        RECT 0.605 1.49 2.735 1.66 ;
        RECT 2.405 1.26 2.735 1.49 ;
    END
    ANTENNAGATEAREA 0.318 LAYER met1 ;
    ANTENNAGATEAREA 0.318 LAYER met2 ;
    ANTENNAGATEAREA 0.318 LAYER met3 ;
    ANTENNAGATEAREA 0.318 LAYER met4 ;
    ANTENNAGATEAREA 0.318 LAYER met5 ;
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.81 2.1 1.265 ;
    END
    ANTENNAGATEAREA 0.159 LAYER met1 ;
    ANTENNAGATEAREA 0.159 LAYER met2 ;
    ANTENNAGATEAREA 0.159 LAYER met3 ;
    ANTENNAGATEAREA 0.159 LAYER met4 ;
    ANTENNAGATEAREA 0.159 LAYER met5 ;
  END D

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.88 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.88 0.245 ;
    END
  END vgnd

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3.935 1.965 10.945 2.105 ;
        RECT 10.655 2.105 10.945 2.15 ;
        RECT 10.655 1.92 10.945 1.965 ;
        RECT 3.935 2.105 4.225 2.15 ;
        RECT 7.775 2.105 8.065 2.15 ;
        RECT 3.935 1.92 4.225 1.965 ;
        RECT 7.775 1.92 8.065 1.965 ;
    END
    ANTENNAGATEAREA 0.411 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.956 LAYER met1 ;
    ANTENNAGATEAREA 0.411 LAYER met2 ;
    ANTENNAGATEAREA 0.411 LAYER met3 ;
    ANTENNAGATEAREA 0.411 LAYER met4 ;
    ANTENNAGATEAREA 0.411 LAYER met5 ;
  END RESETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 1.95 8.005 2.12 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 1.95 4.165 2.12 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 1.95 10.885 2.12 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
    LAYER li1 ;
      RECT 0 3.245 14.88 3.415 ;
      RECT 14.47 2.11 14.765 3.245 ;
      RECT 4.705 2.75 5.035 3.245 ;
      RECT 3.095 2.685 3.425 3.245 ;
      RECT 7.17 2.66 7.52 3.245 ;
      RECT 10.465 2.52 10.795 3.245 ;
      RECT 11.65 1.82 11.9 3.245 ;
      RECT 12.635 1.82 12.885 3.245 ;
      RECT 8.365 1.745 8.535 3.245 ;
      RECT 13.615 2.11 13.865 3.245 ;
      RECT 0.615 2.345 1.565 3.245 ;
      RECT 3.785 1.83 4.165 2.16 ;
      RECT 9.245 2.065 9.955 2.38 ;
      RECT 9.245 1.235 9.415 2.065 ;
      RECT 8.825 0.905 9.415 1.235 ;
      RECT 8.825 0.425 8.995 0.905 ;
      RECT 7.93 0.255 8.995 0.425 ;
      RECT 7.93 0.425 8.1 0.58 ;
      RECT 7.055 0.58 8.1 0.75 ;
      RECT 7.055 0.5 7.225 0.58 ;
      RECT 5.215 0.33 7.225 0.5 ;
      RECT 5.215 0.5 5.62 0.92 ;
      RECT 5.195 0.92 5.62 1.24 ;
      RECT 5.45 1.24 5.62 1.585 ;
      RECT 5.45 1.585 6.205 1.91 ;
      RECT 5.155 1.91 6.205 1.915 ;
      RECT 5.155 1.915 5.655 2.24 ;
      RECT 10.585 1.82 10.915 2.15 ;
      RECT 0 -0.085 14.88 0.085 ;
      RECT 14.435 0.085 14.765 1.13 ;
      RECT 3.67 0.085 3.995 0.75 ;
      RECT 4.715 0.085 5.045 0.75 ;
      RECT 7.43 0.085 7.76 0.41 ;
      RECT 10.14 0.085 10.58 0.68 ;
      RECT 12.105 0.085 12.365 1.1 ;
      RECT 13.035 0.085 13.905 0.76 ;
      RECT 0.545 0.085 0.875 0.765 ;
      RECT 11.755 1.27 13.85 1.6 ;
      RECT 12.1 1.6 12.43 2.7 ;
      RECT 11.755 0.35 11.925 1.27 ;
      RECT 3.615 2.59 3.995 2.98 ;
      RECT 3.615 2.58 4.645 2.59 ;
      RECT 3.615 2.515 6.075 2.58 ;
      RECT 5.745 2.58 6.075 2.755 ;
      RECT 2.105 2.42 6.075 2.515 ;
      RECT 4.58 2.41 6.075 2.42 ;
      RECT 2.105 2.345 3.995 2.42 ;
      RECT 5.825 2.255 6.075 2.41 ;
      RECT 3.445 2.33 3.995 2.345 ;
      RECT 5.825 2.085 6.545 2.255 ;
      RECT 6.375 1.415 6.545 2.085 ;
      RECT 5.79 1.245 6.545 1.415 ;
      RECT 5.79 0.67 5.99 1.245 ;
      RECT 3.445 1.09 3.615 2.33 ;
      RECT 2.565 0.92 3.615 1.09 ;
      RECT 2.105 2.515 2.435 2.98 ;
      RECT 2.565 0.845 2.735 0.92 ;
      RECT 2.27 0.595 2.735 0.845 ;
      RECT 6.245 2.49 6.885 2.755 ;
      RECT 6.245 2.425 8.055 2.49 ;
      RECT 7.725 2.49 8.055 2.755 ;
      RECT 6.715 2.32 8.055 2.425 ;
      RECT 7.495 1.575 7.665 2.32 ;
      RECT 6.715 1.075 6.885 2.32 ;
      RECT 7.495 1.26 8.315 1.575 ;
      RECT 6.16 0.905 6.885 1.075 ;
      RECT 6.16 0.67 6.47 0.905 ;
      RECT 8.735 1.575 9.065 2.755 ;
      RECT 8.485 1.405 9.065 1.575 ;
      RECT 8.485 1.09 8.655 1.405 ;
      RECT 7.055 0.92 8.655 1.09 ;
      RECT 7.055 1.09 7.325 1.945 ;
      RECT 8.27 0.595 8.655 0.92 ;
      RECT 7.835 1.82 8.145 2.15 ;
      RECT 1.105 0.425 1.435 0.64 ;
      RECT 1.105 0.255 3.5 0.425 ;
      RECT 3.225 0.425 3.5 0.75 ;
      RECT 9.27 2.55 10.295 2.88 ;
      RECT 10.125 1.895 10.295 2.55 ;
      RECT 9.585 1.725 10.295 1.895 ;
      RECT 9.585 1.055 9.755 1.725 ;
      RECT 9.585 0.885 11.245 1.055 ;
      RECT 10.915 1.055 11.245 1.215 ;
      RECT 9.585 0.735 9.755 0.885 ;
      RECT 9.165 0.405 9.755 0.735 ;
      RECT 0.115 2.005 2.705 2.175 ;
      RECT 2.375 1.83 2.705 2.005 ;
      RECT 0.115 2.175 0.445 2.98 ;
      RECT 0.115 1.265 0.285 2.005 ;
      RECT 0.115 0.35 0.365 0.935 ;
      RECT 0.115 0.935 1.14 1.265 ;
      RECT 11 2.52 11.33 2.98 ;
      RECT 11.16 1.555 11.33 2.52 ;
      RECT 10.015 1.385 11.585 1.555 ;
      RECT 10.015 1.225 10.345 1.385 ;
      RECT 11.415 0.715 11.585 1.385 ;
      RECT 11.04 0.385 11.585 0.715 ;
      RECT 4.335 1.99 4.515 2.25 ;
      RECT 4.335 1.82 4.975 1.99 ;
      RECT 4.805 1.74 4.975 1.82 ;
      RECT 4.805 1.41 5.28 1.74 ;
      RECT 4.805 1.09 4.975 1.41 ;
      RECT 4.365 0.92 4.975 1.09 ;
      RECT 4.365 0.75 4.535 0.92 ;
      RECT 4.165 0.55 4.535 0.75 ;
  END
END scs8ls_sdfrtp_4

MACRO scs8ls_sdfsbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 14.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.79 1.585 2.12 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.505 1.62 0.835 1.85 ;
        RECT 0.505 1.45 2.045 1.62 ;
        RECT 1.795 1.26 2.045 1.45 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.275 1.18 3.715 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555 1.14 2.765 2.15 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.125 0.35 12.62 1.13 ;
        RECT 12.45 1.13 12.62 1.82 ;
        RECT 12.45 1.82 12.705 2.98 ;
    END
    ANTENNADIFFAREA 0.5357 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.955 0.35 14.29 2.98 ;
    END
    ANTENNADIFFAREA 0.5357 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.4 3.575 ;
    END
  END vpwr

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.295 1.595 9.985 1.735 ;
        RECT 7.295 1.735 7.585 1.78 ;
        RECT 9.695 1.735 9.985 1.78 ;
        RECT 7.295 1.55 7.585 1.595 ;
        RECT 9.695 1.55 9.985 1.595 ;
    END
    ANTENNAGATEAREA 0.252 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.869 LAYER met1 ;
  END SETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.355 1.58 7.525 1.75 ;
      RECT 9.755 1.58 9.925 1.75 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
    LAYER li1 ;
      RECT 6.935 1.915 7.105 2.735 ;
      RECT 6.05 1.69 7.105 1.915 ;
      RECT 2.935 1.99 3.455 2.15 ;
      RECT 2.935 1.82 4.215 1.99 ;
      RECT 3.885 1.22 4.215 1.82 ;
      RECT 2.935 1.01 3.105 1.82 ;
      RECT 2.935 0.34 3.2 1.01 ;
      RECT 5.12 2.37 5.45 2.735 ;
      RECT 5.2 1.52 5.37 2.37 ;
      RECT 5.2 1.35 7.11 1.52 ;
      RECT 6.725 1.19 7.11 1.35 ;
      RECT 5.2 0.35 5.45 1.35 ;
      RECT 6.94 1.075 7.11 1.19 ;
      RECT 6.94 0.905 8.165 1.075 ;
      RECT 7.835 1.075 8.165 1.45 ;
      RECT 4.76 1.37 5.03 2.04 ;
      RECT 4.86 0.425 5.03 1.37 ;
      RECT 3.88 0.255 5.03 0.425 ;
      RECT 3.88 0.425 4.21 1.01 ;
      RECT 5.815 0.905 6.485 1.18 ;
      RECT 5.815 0.735 6.77 0.905 ;
      RECT 6.6 0.35 6.93 0.735 ;
      RECT 13.005 1.55 13.255 2.875 ;
      RECT 13.005 1.22 13.785 1.55 ;
      RECT 13.005 1.13 13.255 1.22 ;
      RECT 12.84 0.54 13.255 1.13 ;
      RECT 2.215 2.38 3.795 2.49 ;
      RECT 2.215 2.32 4.925 2.38 ;
      RECT 4.59 2.38 4.925 2.735 ;
      RECT 3.625 2.21 4.925 2.32 ;
      RECT 4.42 0.925 4.59 2.21 ;
      RECT 4.42 0.595 4.69 0.925 ;
      RECT 1.435 2.8 1.945 2.96 ;
      RECT 1.435 2.63 2.385 2.8 ;
      RECT 2.215 2.49 2.385 2.63 ;
      RECT 2.215 1.09 2.385 2.32 ;
      RECT 1.505 0.92 2.385 1.09 ;
      RECT 1.505 0.35 1.835 0.92 ;
      RECT 7.985 2.52 8.315 2.755 ;
      RECT 7.985 2.35 9.83 2.52 ;
      RECT 9.58 2.52 9.83 2.735 ;
      RECT 7.985 2.29 8.315 2.35 ;
      RECT 9.58 2.29 9.83 2.35 ;
      RECT 8.53 2.905 10.38 3.075 ;
      RECT 8.53 2.69 8.86 2.905 ;
      RECT 10.05 2.52 10.38 2.905 ;
      RECT 10.95 2.52 11.28 2.98 ;
      RECT 11.11 2.265 11.28 2.52 ;
      RECT 10 2.12 11.28 2.265 ;
      RECT 9.045 2.095 11.28 2.12 ;
      RECT 9.045 2.12 9.38 2.18 ;
      RECT 11.11 1.97 11.28 2.095 ;
      RECT 9.045 1.95 10.17 2.095 ;
      RECT 11.11 1.64 11.895 1.97 ;
      RECT 9.045 1.85 9.38 1.95 ;
      RECT 9.21 1.05 9.38 1.85 ;
      RECT 8.785 0.35 9.38 1.05 ;
      RECT 11.5 2.18 12.235 2.35 ;
      RECT 12.065 1.47 12.235 2.18 ;
      RECT 11.225 1.3 12.235 1.47 ;
      RECT 11.5 2.35 11.75 2.98 ;
      RECT 11.225 1.07 11.395 1.3 ;
      RECT 9.62 0.9 11.395 1.07 ;
      RECT 9.62 1.07 9.95 1.23 ;
      RECT 11.065 0.35 11.395 0.9 ;
      RECT 4.105 2.905 5.81 3.075 ;
      RECT 4.105 2.55 4.355 2.905 ;
      RECT 5.64 2.255 5.81 2.905 ;
      RECT 5.64 2.085 6.765 2.255 ;
      RECT 6.595 2.255 6.765 2.905 ;
      RECT 5.64 2.02 5.81 2.085 ;
      RECT 6.595 2.905 7.445 3.075 ;
      RECT 5.54 1.69 5.81 2.02 ;
      RECT 7.275 2.12 7.445 2.905 ;
      RECT 7.275 1.95 8.83 2.12 ;
      RECT 8.66 1.68 8.83 1.95 ;
      RECT 8.66 1.35 8.99 1.68 ;
      RECT 7.295 1.245 7.625 1.78 ;
      RECT 0.115 2.29 2.045 2.46 ;
      RECT 1.795 1.83 2.045 2.29 ;
      RECT 0.115 2.46 0.365 2.98 ;
      RECT 0.115 1.28 0.335 2.29 ;
      RECT 0.115 0.35 0.445 0.95 ;
      RECT 0.115 0.95 1.14 1.28 ;
      RECT 10.585 1.78 10.915 1.925 ;
      RECT 9.725 1.55 10.915 1.78 ;
      RECT 10.585 1.255 10.915 1.55 ;
      RECT 0 3.245 14.4 3.415 ;
      RECT 13.455 1.995 13.785 3.245 ;
      RECT 2.555 2.66 2.82 3.245 ;
      RECT 3.575 2.66 3.905 3.245 ;
      RECT 10.58 2.52 10.75 3.245 ;
      RECT 11.95 2.52 12.28 3.245 ;
      RECT 6.175 2.425 6.425 3.245 ;
      RECT 7.615 2.295 7.785 3.245 ;
      RECT 0.565 2.63 0.895 3.245 ;
      RECT 0 -0.085 14.4 0.085 ;
      RECT 13.455 0.085 13.785 1.05 ;
      RECT 0.615 0.085 0.945 0.78 ;
      RECT 2.325 0.085 2.655 0.75 ;
      RECT 3.38 0.085 3.71 1.01 ;
      RECT 6.02 0.085 6.37 0.565 ;
      RECT 7.5 0.085 8.295 0.735 ;
      RECT 10.285 0.085 10.895 0.68 ;
      RECT 11.625 0.085 11.955 1.13 ;
  END
END scs8ls_sdfsbp_1

MACRO scs8ls_sdfsbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 17.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965 0.9 2.295 1.4 ;
        RECT 0.425 1.4 2.295 1.57 ;
        RECT 0.425 1.57 1.085 1.8 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.385 0.44 1.795 1.23 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.715 1.18 4.195 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.885 0.35 17.225 1.13 ;
        RECT 17.055 1.13 17.225 1.82 ;
        RECT 16.865 1.82 17.225 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.85 0.35 15.235 1.41 ;
        RECT 14.85 1.41 15.105 2.98 ;
    END
    ANTENNADIFFAREA 0.558 ;
  END QN

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.805 0.95 3.205 1.62 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 17.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 17.76 3.575 ;
    END
  END vpwr

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.775 1.595 13.345 1.735 ;
        RECT 13.055 1.735 13.345 1.78 ;
        RECT 13.055 1.55 13.345 1.595 ;
        RECT 7.775 1.735 8.065 1.78 ;
        RECT 7.775 1.55 8.065 1.595 ;
    END
    ANTENNAGATEAREA 0.252 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 3.885 LAYER met1 ;
  END SETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.835 1.58 8.005 1.75 ;
      RECT 13.115 1.58 13.285 1.75 ;
      RECT 17.435 -0.085 17.605 0.085 ;
      RECT 16.955 -0.085 17.125 0.085 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 17.435 3.245 17.605 3.415 ;
      RECT 16.955 3.245 17.125 3.415 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
    LAYER li1 ;
      RECT 6.815 1.04 7.145 1.225 ;
      RECT 6.815 0.87 7.71 1.04 ;
      RECT 7.38 0.35 7.71 0.87 ;
      RECT 7.495 2.295 7.825 2.735 ;
      RECT 7.495 1.995 7.665 2.295 ;
      RECT 6.635 1.735 7.665 1.995 ;
      RECT 8.735 1.87 9.065 1.96 ;
      RECT 8.735 1.7 12.05 1.87 ;
      RECT 8.735 1.685 9.065 1.7 ;
      RECT 11.72 0.9 12.05 1.7 ;
      RECT 3.075 1.79 4.72 1.96 ;
      RECT 4.39 1.35 4.72 1.79 ;
      RECT 3.075 1.96 3.545 2.14 ;
      RECT 3.375 1.01 3.545 1.79 ;
      RECT 3.375 0.34 3.65 1.01 ;
      RECT 4.39 2.905 6.24 3.075 ;
      RECT 4.39 2.47 4.72 2.905 ;
      RECT 6.07 2.335 6.24 2.905 ;
      RECT 6.07 2.165 7.325 2.335 ;
      RECT 7.155 2.335 7.325 2.905 ;
      RECT 6.07 0.97 6.305 2.165 ;
      RECT 7.155 2.905 8.165 3.075 ;
      RECT 7.995 2.22 8.165 2.905 ;
      RECT 7.995 2.05 8.565 2.22 ;
      RECT 8.395 1.515 8.565 2.05 ;
      RECT 8.395 1.345 11.39 1.515 ;
      RECT 10.38 1.515 11.39 1.53 ;
      RECT 10.38 1.2 11.39 1.345 ;
      RECT 5.23 1.29 5.56 1.96 ;
      RECT 5.39 0.425 5.56 1.29 ;
      RECT 4.33 0.255 5.56 0.425 ;
      RECT 4.33 0.425 4.66 1.01 ;
      RECT 9.03 1.005 10.21 1.175 ;
      RECT 9.96 0.425 10.21 1.005 ;
      RECT 9.03 0.35 9.28 1.005 ;
      RECT 9.96 0.255 11.21 0.425 ;
      RECT 10.88 0.425 11.21 0.69 ;
      RECT 1.505 2.31 3.885 2.48 ;
      RECT 3.715 2.3 3.885 2.31 ;
      RECT 3.715 2.13 5.37 2.3 ;
      RECT 4.89 2.3 5.37 2.735 ;
      RECT 4.89 0.845 5.06 2.13 ;
      RECT 4.89 0.595 5.22 0.845 ;
      RECT 2.465 0.73 2.635 2.31 ;
      RECT 1.965 0.56 2.635 0.73 ;
      RECT 1.965 0.4 2.35 0.56 ;
      RECT 1.505 2.48 1.955 2.98 ;
      RECT 5.54 2.295 5.9 2.735 ;
      RECT 5.73 0.8 5.9 2.295 ;
      RECT 5.73 0.47 6.645 0.8 ;
      RECT 6.475 0.8 6.645 1.395 ;
      RECT 6.475 1.395 7.665 1.565 ;
      RECT 7.355 1.38 7.665 1.395 ;
      RECT 7.355 1.21 8.05 1.38 ;
      RECT 7.88 1.175 8.05 1.21 ;
      RECT 7.88 0.9 8.86 1.175 ;
      RECT 9.875 2.905 11.105 3.075 ;
      RECT 10.775 2.38 11.105 2.905 ;
      RECT 9.875 2.3 10.125 2.905 ;
      RECT 8.925 2.13 10.125 2.3 ;
      RECT 8.925 2.3 9.255 2.98 ;
      RECT 9.875 2.1 10.125 2.13 ;
      RECT 11.365 2.885 12.74 3.055 ;
      RECT 12.41 2.52 12.74 2.885 ;
      RECT 11.365 2.385 11.62 2.885 ;
      RECT 11.82 2.31 12.22 2.715 ;
      RECT 11.82 2.21 13.975 2.31 ;
      RECT 13.31 2.31 13.64 2.98 ;
      RECT 10.325 2.14 13.975 2.21 ;
      RECT 10.325 2.21 10.575 2.7 ;
      RECT 10.325 2.04 12.39 2.14 ;
      RECT 13.645 1.3 13.975 2.14 ;
      RECT 12.22 0.73 12.39 2.04 ;
      RECT 11.38 0.4 12.39 0.73 ;
      RECT 11.38 0.73 11.55 0.86 ;
      RECT 10.38 0.86 11.55 1.03 ;
      RECT 10.38 0.595 10.71 0.86 ;
      RECT 13.87 2.48 14.315 2.91 ;
      RECT 14.145 1.13 14.315 2.48 ;
      RECT 12.565 0.96 14.315 1.13 ;
      RECT 12.565 1.13 12.895 1.96 ;
      RECT 13.77 0.35 14.1 0.96 ;
      RECT 15.865 1.3 16.885 1.63 ;
      RECT 15.865 1.63 16.195 2.86 ;
      RECT 15.865 0.45 16.22 1.3 ;
      RECT 7.835 1.55 8.225 1.88 ;
      RECT 0.085 1.97 2.105 2.14 ;
      RECT 1.775 1.81 2.105 1.97 ;
      RECT 0.085 1.23 0.255 1.97 ;
      RECT 0.085 2.14 0.465 2.98 ;
      RECT 0.085 0.9 1.145 1.23 ;
      RECT 0.085 0.35 0.445 0.9 ;
      RECT 13.085 1.3 13.435 1.97 ;
      RECT 0 -0.085 17.76 0.085 ;
      RECT 17.395 0.085 17.645 1.13 ;
      RECT 15.405 0.085 15.655 1.13 ;
      RECT 16.455 0.085 16.705 1.13 ;
      RECT 2.84 0.085 3.17 0.78 ;
      RECT 3.83 0.085 4.16 1.01 ;
      RECT 6.815 0.085 7.15 0.7 ;
      RECT 8.2 0.085 8.53 0.68 ;
      RECT 9.45 0.085 9.78 0.835 ;
      RECT 13.26 0.085 13.59 0.79 ;
      RECT 14.35 0.085 14.68 0.79 ;
      RECT 0.615 0.085 1.02 0.68 ;
      RECT 0 3.245 17.76 3.415 ;
      RECT 17.395 1.82 17.645 3.245 ;
      RECT 15.305 1.82 15.635 3.245 ;
      RECT 16.415 1.82 16.665 3.245 ;
      RECT 2.495 2.65 2.845 3.245 ;
      RECT 3.525 2.65 4.22 3.245 ;
      RECT 12.94 2.52 13.11 3.245 ;
      RECT 6.41 2.505 6.985 3.245 ;
      RECT 9.425 2.47 9.675 3.245 ;
      RECT 8.335 2.39 8.665 3.245 ;
      RECT 0.635 2.31 0.965 3.245 ;
      RECT 14.485 1.82 14.655 3.245 ;
  END
END scs8ls_sdfsbp_2

MACRO scs8ls_sdfstp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 13.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.82 1.58 2.15 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.61 0.835 1.95 ;
        RECT 0.425 1.44 2.045 1.61 ;
        RECT 0.425 1.28 0.68 1.44 ;
        RECT 1.79 1.26 2.045 1.44 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.315 1.18 3.715 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555 1.14 2.805 2.15 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.38 0.35 13.815 1.05 ;
        RECT 13.565 1.05 13.815 2.98 ;
    END
    ANTENNADIFFAREA 0.5301 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.92 3.575 ;
    END
  END vpwr

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.295 1.595 10.945 1.735 ;
        RECT 7.295 1.735 7.585 1.78 ;
        RECT 10.655 1.735 10.945 1.78 ;
        RECT 7.295 1.55 7.585 1.595 ;
        RECT 10.655 1.55 10.945 1.595 ;
    END
    ANTENNAGATEAREA 0.252 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.541 LAYER met1 ;
  END SETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.355 1.58 7.525 1.75 ;
      RECT 10.715 1.58 10.885 1.75 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
    LAYER li1 ;
      RECT 4.785 1.105 5.005 2.07 ;
      RECT 4.785 0.935 5.205 1.105 ;
      RECT 5.035 0.425 5.205 0.935 ;
      RECT 3.975 0.255 5.205 0.425 ;
      RECT 3.975 0.425 4.225 1.13 ;
      RECT 2.975 1.82 4.215 2.07 ;
      RECT 3.885 1.35 4.215 1.82 ;
      RECT 2.975 1.01 3.145 1.82 ;
      RECT 2.975 0.35 3.305 1.01 ;
      RECT 4.105 2.895 5.845 3.065 ;
      RECT 4.105 2.58 4.275 2.895 ;
      RECT 5.675 2.515 5.845 2.895 ;
      RECT 5.675 2.345 6.815 2.515 ;
      RECT 6.645 2.515 6.815 2.895 ;
      RECT 5.675 1.945 5.845 2.345 ;
      RECT 6.645 2.895 7.495 3.065 ;
      RECT 5.515 1.775 5.845 1.945 ;
      RECT 7.325 2.14 7.495 2.895 ;
      RECT 5.515 1.615 5.73 1.775 ;
      RECT 7.325 1.97 7.945 2.14 ;
      RECT 7.775 1.75 7.945 1.97 ;
      RECT 7.775 1.58 8.84 1.75 ;
      RECT 8.67 1.45 8.84 1.58 ;
      RECT 8.67 1.12 9 1.45 ;
      RECT 6.24 1.03 6.48 1.265 ;
      RECT 6.24 0.86 7.005 1.03 ;
      RECT 6.675 0.57 7.005 0.86 ;
      RECT 12.53 1.22 13.395 1.55 ;
      RECT 12.53 1.995 12.86 2.875 ;
      RECT 12.53 1.55 12.7 1.995 ;
      RECT 12.53 1.005 12.7 1.22 ;
      RECT 12.37 0.87 12.7 1.005 ;
      RECT 11.955 0.54 12.7 0.87 ;
      RECT 2.215 2.49 3.405 2.66 ;
      RECT 3.235 2.41 3.405 2.49 ;
      RECT 3.235 2.24 5.005 2.41 ;
      RECT 4.445 2.41 5.005 2.725 ;
      RECT 4.445 0.765 4.615 2.24 ;
      RECT 4.445 0.595 4.865 0.765 ;
      RECT 1.43 2.66 2.385 2.91 ;
      RECT 2.215 1.09 2.385 2.49 ;
      RECT 1.555 0.92 2.385 1.09 ;
      RECT 1.555 0.35 1.885 0.92 ;
      RECT 5.175 2.265 5.505 2.725 ;
      RECT 5.175 1.445 5.345 2.265 ;
      RECT 5.175 1.435 6.935 1.445 ;
      RECT 5.9 1.445 6.935 1.605 ;
      RECT 6.65 1.37 6.935 1.435 ;
      RECT 5.175 1.275 6.07 1.435 ;
      RECT 6.65 1.605 6.935 1.835 ;
      RECT 6.65 1.2 8.43 1.37 ;
      RECT 5.375 0.385 5.625 1.275 ;
      RECT 7.76 1.37 8.43 1.41 ;
      RECT 7.76 1.12 8.43 1.2 ;
      RECT 8.115 2.52 8.365 2.725 ;
      RECT 8.115 2.35 9.895 2.52 ;
      RECT 9.565 2.52 9.895 2.735 ;
      RECT 9.565 1.96 9.895 2.35 ;
      RECT 8.115 1.92 8.365 2.35 ;
      RECT 8.585 2.905 10.43 3.075 ;
      RECT 8.585 2.69 8.915 2.905 ;
      RECT 10.1 2.56 10.43 2.905 ;
      RECT 11 2.39 11.37 2.98 ;
      RECT 10.065 2.22 11.37 2.39 ;
      RECT 11.2 2.05 11.37 2.22 ;
      RECT 10.065 1.79 10.235 2.22 ;
      RECT 11.2 1.38 11.6 2.05 ;
      RECT 9.09 1.62 10.235 1.79 ;
      RECT 9.09 1.79 9.365 2.18 ;
      RECT 9.195 0.94 9.365 1.62 ;
      RECT 8.795 0.35 9.365 0.94 ;
      RECT 11.54 2.39 11.87 2.98 ;
      RECT 11.54 2.22 11.94 2.39 ;
      RECT 11.77 1.21 11.94 2.22 ;
      RECT 9.79 1.04 11.94 1.21 ;
      RECT 9.79 1.21 10.46 1.31 ;
      RECT 9.79 0.98 11.77 1.04 ;
      RECT 11.395 0.35 11.77 0.98 ;
      RECT 7.145 1.54 7.555 1.8 ;
      RECT 0.085 2.32 2.045 2.49 ;
      RECT 1.79 1.83 2.045 2.32 ;
      RECT 0.085 2.49 0.36 2.98 ;
      RECT 0.085 2.3 0.36 2.32 ;
      RECT 0.085 1.11 0.255 2.3 ;
      RECT 0.085 0.94 1.22 1.11 ;
      RECT 0.89 1.11 1.22 1.27 ;
      RECT 0.085 0.35 0.525 0.94 ;
      RECT 10.685 1.38 11.03 2.05 ;
      RECT 0 3.245 13.92 3.415 ;
      RECT 2.565 2.83 2.895 3.245 ;
      RECT 6.225 2.685 6.475 3.245 ;
      RECT 3.575 2.58 3.905 3.245 ;
      RECT 10.63 2.56 10.8 3.245 ;
      RECT 12.07 2.56 12.32 3.245 ;
      RECT 7.665 2.31 7.915 3.245 ;
      RECT 13.03 1.995 13.36 3.245 ;
      RECT 0.56 2.66 0.89 3.245 ;
      RECT 0 -0.085 13.92 0.085 ;
      RECT 0.695 0.085 1.025 0.77 ;
      RECT 2.375 0.085 2.705 0.75 ;
      RECT 3.475 0.085 3.805 1.01 ;
      RECT 6.115 0.085 6.445 0.69 ;
      RECT 7.455 0.085 8.305 0.94 ;
      RECT 10.825 0.085 11.155 0.81 ;
      RECT 12.88 0.085 13.21 1.05 ;
      RECT 6.985 2.175 7.155 2.725 ;
      RECT 6.015 2.005 7.155 2.175 ;
      RECT 6.015 1.795 6.345 2.005 ;
  END
END scs8ls_sdfstp_1

MACRO scs8ls_sdfstp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 14.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.325 1.49 14.755 1.82 ;
        RECT 13.995 1.82 14.755 2.15 ;
        RECT 14.175 1.32 14.755 1.49 ;
        RECT 13.995 2.15 14.275 2.98 ;
        RECT 14.175 1.15 14.345 1.32 ;
        RECT 13.99 0.37 14.345 1.15 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END Q

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555 1.14 2.78 2.15 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.82 1.585 2.15 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475 1.58 0.805 2.14 ;
        RECT 0.475 1.41 2.045 1.58 ;
        RECT 1.795 1.25 2.045 1.41 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.3 1.18 3.715 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.88 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.88 0.245 ;
    END
  END vgnd

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.295 1.225 11.905 1.365 ;
        RECT 7.295 1.365 7.585 1.41 ;
        RECT 11.615 1.365 11.905 1.41 ;
        RECT 7.295 1.18 7.585 1.225 ;
        RECT 11.615 1.18 11.905 1.225 ;
    END
    ANTENNAGATEAREA 0.252 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 3.213 LAYER met1 ;
  END SETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.355 1.21 7.525 1.38 ;
      RECT 11.675 1.21 11.845 1.38 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
    LAYER li1 ;
      RECT 8.18 0.885 10.08 1.055 ;
      RECT 9.75 0.595 10.08 0.885 ;
      RECT 8.18 0.35 8.51 0.885 ;
      RECT 7.905 2.235 8.235 2.755 ;
      RECT 7.905 2.145 8.765 2.235 ;
      RECT 7.905 2.065 9.83 2.145 ;
      RECT 9.5 2.145 9.83 2.735 ;
      RECT 8.595 1.975 9.83 2.065 ;
      RECT 6.515 2.905 7.365 3.075 ;
      RECT 6.515 2.255 6.685 2.905 ;
      RECT 7.195 1.895 7.365 2.905 ;
      RECT 5.56 2.085 6.685 2.255 ;
      RECT 7.195 1.805 8.425 1.895 ;
      RECT 5.56 2.255 5.73 2.895 ;
      RECT 5.56 2.045 5.73 2.085 ;
      RECT 7.195 1.725 10.17 1.805 ;
      RECT 4.075 2.895 5.73 3.065 ;
      RECT 5.475 1.715 5.73 2.045 ;
      RECT 10 1.805 10.72 2.135 ;
      RECT 8.255 1.475 10.17 1.725 ;
      RECT 4.075 2.58 4.325 2.895 ;
      RECT 5.98 0.7 6.31 1.205 ;
      RECT 5.98 0.53 7.02 0.7 ;
      RECT 6.69 0.35 7.02 0.53 ;
      RECT 6.855 1.915 7.025 2.735 ;
      RECT 5.94 1.745 7.025 1.915 ;
      RECT 5.94 1.715 6.27 1.745 ;
      RECT 2.96 1.82 4.215 2.07 ;
      RECT 3.885 1.35 4.215 1.82 ;
      RECT 2.96 0.35 3.35 1.01 ;
      RECT 2.96 1.01 3.13 1.82 ;
      RECT 5.115 2.265 5.365 2.725 ;
      RECT 5.135 1.545 5.305 2.265 ;
      RECT 5.135 1.375 6.88 1.545 ;
      RECT 6.55 1.545 6.88 1.57 ;
      RECT 6.55 1.04 6.88 1.375 ;
      RECT 5.34 0.385 5.59 1.375 ;
      RECT 6.55 0.87 7.925 1.04 ;
      RECT 7.755 1.04 7.925 1.225 ;
      RECT 7.755 1.225 8.085 1.555 ;
      RECT 4.76 1.185 4.965 1.73 ;
      RECT 4.76 1.015 5.17 1.185 ;
      RECT 5 0.425 5.17 1.015 ;
      RECT 4.03 0.255 5.17 0.425 ;
      RECT 4.03 0.425 4.2 1.13 ;
      RECT 13.035 1.32 14.005 1.65 ;
      RECT 13.035 1.65 13.37 2.98 ;
      RECT 13.035 0.47 13.365 1.32 ;
      RECT 9 2.905 10.435 3.075 ;
      RECT 10.105 2.475 10.435 2.905 ;
      RECT 9 2.315 9.33 2.905 ;
      RECT 10.105 2.305 11.86 2.475 ;
      RECT 11.53 2.475 11.86 2.98 ;
      RECT 10.89 2.14 11.86 2.305 ;
      RECT 10.89 1.97 12.465 2.14 ;
      RECT 10.89 1.57 11.06 1.97 ;
      RECT 12.135 1.13 12.465 1.97 ;
      RECT 10.41 1.4 11.06 1.57 ;
      RECT 10.41 0.81 10.58 1.4 ;
      RECT 10.25 0.425 10.58 0.81 ;
      RECT 9.25 0.255 10.58 0.425 ;
      RECT 9.25 0.425 9.58 0.715 ;
      RECT 7.205 1.21 7.555 1.555 ;
      RECT 2.95 2.24 4.915 2.41 ;
      RECT 4.585 2.41 4.915 2.725 ;
      RECT 4.585 2.07 4.915 2.24 ;
      RECT 4.42 1.9 4.915 2.07 ;
      RECT 4.42 0.845 4.59 1.9 ;
      RECT 4.42 0.595 4.83 0.845 ;
      RECT 2.215 2.49 3.12 2.66 ;
      RECT 2.95 2.41 3.12 2.49 ;
      RECT 1.435 2.66 2.385 2.91 ;
      RECT 2.215 1.08 2.385 2.49 ;
      RECT 1.56 0.91 2.385 1.08 ;
      RECT 1.56 0.35 1.89 0.91 ;
      RECT 11.445 1.18 11.875 1.8 ;
      RECT 12.06 2.48 12.31 2.98 ;
      RECT 12.06 2.31 12.805 2.48 ;
      RECT 12.635 0.96 12.805 2.31 ;
      RECT 10.945 0.79 12.805 0.96 ;
      RECT 10.945 0.96 11.275 1.23 ;
      RECT 12.5 0.35 12.805 0.79 ;
      RECT 0 -0.085 14.88 0.085 ;
      RECT 14.515 0.085 14.765 1.15 ;
      RECT 2.46 0.085 2.79 0.74 ;
      RECT 3.52 0.085 3.85 1.01 ;
      RECT 6.13 0.085 6.46 0.36 ;
      RECT 7.51 0.085 8.01 0.68 ;
      RECT 8.69 0.085 9.02 0.715 ;
      RECT 11.64 0.085 12.33 0.6 ;
      RECT 13.555 0.085 13.805 1.15 ;
      RECT 0.615 0.085 1.07 0.68 ;
      RECT 0 3.245 14.88 3.415 ;
      RECT 14.445 2.32 14.775 3.245 ;
      RECT 2.56 2.83 2.89 3.245 ;
      RECT 12.51 2.65 12.84 3.245 ;
      RECT 11.08 2.645 11.33 3.245 ;
      RECT 3.545 2.58 3.875 3.245 ;
      RECT 6.095 2.425 6.345 3.245 ;
      RECT 8.435 2.405 8.685 3.245 ;
      RECT 7.535 2.065 7.705 3.245 ;
      RECT 13.54 1.82 13.825 3.245 ;
      RECT 0.565 2.66 0.895 3.245 ;
      RECT 0.115 2.32 2.045 2.49 ;
      RECT 1.795 1.83 2.045 2.32 ;
      RECT 0.115 2.49 0.365 2.98 ;
      RECT 0.115 2.31 0.365 2.32 ;
      RECT 0.115 1.23 0.285 2.31 ;
      RECT 0.115 0.35 0.445 0.9 ;
      RECT 0.115 0.9 1.225 1.23 ;
  END
END scs8ls_sdfstp_2

MACRO scs8ls_sdfstp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 15.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.025 1.61 15.715 1.78 ;
        RECT 15.025 1.78 15.195 1.82 ;
        RECT 15.485 1.44 15.715 1.61 ;
        RECT 14.045 1.82 15.195 2.15 ;
        RECT 14.895 1.27 15.715 1.44 ;
        RECT 14.045 2.15 14.325 2.98 ;
        RECT 15.025 2.15 15.195 2.98 ;
        RECT 14.895 1.15 15.225 1.27 ;
        RECT 13.895 0.98 15.225 1.15 ;
        RECT 13.895 0.35 14.225 0.98 ;
        RECT 14.895 0.35 15.225 0.98 ;
    END
    ANTENNADIFFAREA 1.2011 ;
  END Q

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555 1.1 2.835 2.15 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.105 1.82 1.575 2.15 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.58 0.855 2.15 ;
        RECT 0.525 1.41 2.045 1.58 ;
        RECT 1.715 1.25 2.045 1.41 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.345 1.18 3.715 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 15.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 15.84 3.575 ;
    END
  END vpwr

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.295 1.595 11.905 1.735 ;
        RECT 7.295 1.735 7.585 1.78 ;
        RECT 11.615 1.735 11.905 1.78 ;
        RECT 7.295 1.55 7.585 1.595 ;
        RECT 11.615 1.55 11.905 1.595 ;
    END
    ANTENNAGATEAREA 0.252 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 3.213 LAYER met1 ;
  END SETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.355 1.58 7.525 1.75 ;
      RECT 11.675 1.58 11.845 1.75 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 13.595 -0.085 13.765 0.085 ;
    LAYER li1 ;
      RECT 10.545 2.65 10.955 2.98 ;
      RECT 13.17 1.49 14.695 1.65 ;
      RECT 12.88 1.32 14.695 1.49 ;
      RECT 13.17 1.65 13.34 2.98 ;
      RECT 12.88 0.35 13.21 1.32 ;
      RECT 8.085 2.29 8.365 2.715 ;
      RECT 8.085 2.12 9.875 2.29 ;
      RECT 9.545 2.29 9.875 2.69 ;
      RECT 9.545 2.1 9.875 2.12 ;
      RECT 4.07 2.895 5.83 3.065 ;
      RECT 4.07 2.58 4.4 2.895 ;
      RECT 5.66 2.46 5.83 2.895 ;
      RECT 5.66 2.29 6.865 2.46 ;
      RECT 6.695 2.46 6.865 2.895 ;
      RECT 5.66 2.105 5.83 2.29 ;
      RECT 6.695 2.895 7.545 3.065 ;
      RECT 5.54 1.775 5.83 2.105 ;
      RECT 7.375 2.12 7.545 2.895 ;
      RECT 7.375 1.95 7.895 2.12 ;
      RECT 7.725 1.93 9.375 1.95 ;
      RECT 7.725 1.78 10.765 1.93 ;
      RECT 10.435 1.93 10.765 2.135 ;
      RECT 9.045 1.76 10.765 1.78 ;
      RECT 9.045 1.45 9.375 1.76 ;
      RECT 6.005 0.94 6.335 1.265 ;
      RECT 6.005 0.77 7.1 0.94 ;
      RECT 6.77 0.35 7.1 0.77 ;
      RECT 9.095 2.86 10.375 3.075 ;
      RECT 9.095 2.6 9.375 2.86 ;
      RECT 10.045 2.48 10.375 2.86 ;
      RECT 10.045 2.31 12.21 2.48 ;
      RECT 11.575 2.48 11.905 2.98 ;
      RECT 12.04 2.01 12.21 2.31 ;
      RECT 10.935 1.57 11.105 2.31 ;
      RECT 12.04 1.34 12.37 2.01 ;
      RECT 10.21 1.4 11.105 1.57 ;
      RECT 10.21 0.425 10.54 1.4 ;
      RECT 9.35 0.255 10.54 0.425 ;
      RECT 9.35 0.425 9.68 0.94 ;
      RECT 7.035 2.12 7.205 2.725 ;
      RECT 6.04 1.95 7.205 2.12 ;
      RECT 6.04 1.78 6.37 1.95 ;
      RECT 3.005 1.82 4.215 2.07 ;
      RECT 3.885 1.35 4.215 1.82 ;
      RECT 3.005 0.35 3.39 1.01 ;
      RECT 3.005 1.01 3.175 1.82 ;
      RECT 5.2 2.275 5.48 2.725 ;
      RECT 5.2 1.605 5.37 2.275 ;
      RECT 5.2 1.435 6.955 1.605 ;
      RECT 6.625 1.605 6.955 1.78 ;
      RECT 6.625 1.28 6.955 1.435 ;
      RECT 5.31 0.385 5.64 1.435 ;
      RECT 6.625 1.11 8.265 1.28 ;
      RECT 7.935 1.28 8.265 1.45 ;
      RECT 4.75 1.265 5.03 1.73 ;
      RECT 4.75 1.095 5.14 1.265 ;
      RECT 4.97 0.425 5.14 1.095 ;
      RECT 4.07 0.255 5.14 0.425 ;
      RECT 4.07 0.425 4.24 1.13 ;
      RECT 8.44 1.11 10.03 1.28 ;
      RECT 9.86 0.595 10.03 1.11 ;
      RECT 8.44 0.35 8.61 1.11 ;
      RECT 7.195 1.45 7.555 1.78 ;
      RECT 3.005 2.24 5.03 2.41 ;
      RECT 4.7 2.41 5.03 2.725 ;
      RECT 4.41 1.9 5.03 2.24 ;
      RECT 4.41 0.925 4.58 1.9 ;
      RECT 4.41 0.595 4.8 0.925 ;
      RECT 2.215 2.49 3.175 2.66 ;
      RECT 3.005 2.41 3.175 2.49 ;
      RECT 1.425 2.66 2.385 2.91 ;
      RECT 2.215 1.08 2.385 2.49 ;
      RECT 1.79 0.91 2.385 1.08 ;
      RECT 1.79 0.74 1.96 0.91 ;
      RECT 1.475 0.41 1.96 0.74 ;
      RECT 11.47 1.47 11.87 2.14 ;
      RECT 12.135 2.65 12.55 2.98 ;
      RECT 12.38 2.35 12.55 2.65 ;
      RECT 12.38 2.18 12.71 2.35 ;
      RECT 12.54 1.07 12.71 2.18 ;
      RECT 10.955 0.9 12.71 1.07 ;
      RECT 10.955 1.07 11.285 1.23 ;
      RECT 12.32 0.35 12.71 0.9 ;
      RECT 0 -0.085 15.84 0.085 ;
      RECT 15.395 0.085 15.725 1.1 ;
      RECT 2.45 0.085 2.78 0.74 ;
      RECT 3.56 0.085 3.89 1.01 ;
      RECT 6.21 0.085 6.54 0.6 ;
      RECT 7.59 0.085 8.26 0.93 ;
      RECT 8.79 0.085 9.12 0.94 ;
      RECT 11.65 0.085 12.15 0.68 ;
      RECT 13.38 0.085 13.71 1.13 ;
      RECT 14.395 0.085 14.725 0.81 ;
      RECT 0.615 0.085 0.945 0.74 ;
      RECT 0 3.245 15.84 3.415 ;
      RECT 15.395 1.95 15.725 3.245 ;
      RECT 2.56 2.83 2.89 3.245 ;
      RECT 11.125 2.65 11.375 3.245 ;
      RECT 6.275 2.63 6.525 3.245 ;
      RECT 3.57 2.58 3.9 3.245 ;
      RECT 12.72 2.52 12.97 3.245 ;
      RECT 8.535 2.46 8.865 3.245 ;
      RECT 7.715 2.29 7.885 3.245 ;
      RECT 13.54 2.1 13.87 3.245 ;
      RECT 14.495 2.32 14.825 3.245 ;
      RECT 0.555 2.66 0.885 3.245 ;
      RECT 0.105 2.32 2.045 2.49 ;
      RECT 1.785 1.83 2.045 2.32 ;
      RECT 0.105 2.49 0.355 2.98 ;
      RECT 0.105 1.24 0.355 2.32 ;
      RECT 0.105 0.35 0.445 0.91 ;
      RECT 0.105 0.91 1.14 1.24 ;
  END
END scs8ls_sdfstp_4

MACRO scs8ls_sdfxbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.48 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.38 1.55 2.725 2.15 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.81 2.05 0.955 ;
        RECT 0.425 0.955 2.05 1.285 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.455 1.63 1.785 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.235 1.18 3.685 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.5 0.35 10.915 1.13 ;
        RECT 10.745 1.13 10.915 1.82 ;
        RECT 10.65 1.82 10.915 2.98 ;
    END
    ANTENNADIFFAREA 0.5189 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.035 0.35 12.375 1.05 ;
        RECT 12.155 1.05 12.375 1.82 ;
        RECT 12.045 1.82 12.375 2.98 ;
    END
    ANTENNADIFFAREA 0.5301 ;
  END QN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12.48 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12.48 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
    LAYER li1 ;
      RECT 5.41 2.46 5.765 2.92 ;
      RECT 5.41 1.7 5.58 2.46 ;
      RECT 5.41 1.53 7.02 1.7 ;
      RECT 6.69 1.7 7.02 1.93 ;
      RECT 5.41 0.595 5.58 1.53 ;
      RECT 9.78 1.32 10.575 1.65 ;
      RECT 9.6 2.35 9.95 2.98 ;
      RECT 8.71 2.12 9.95 2.35 ;
      RECT 9.6 1.94 9.95 2.12 ;
      RECT 9.78 1.65 9.95 1.94 ;
      RECT 9.78 0.93 9.95 1.32 ;
      RECT 9.59 0.35 9.95 0.93 ;
      RECT 6.985 2.1 7.395 2.35 ;
      RECT 7.19 1.36 7.36 2.1 ;
      RECT 6.245 1.03 7.36 1.36 ;
      RECT 7.19 0.92 7.36 1.03 ;
      RECT 7.19 0.595 7.52 0.92 ;
      RECT 11.09 1.55 11.34 2.875 ;
      RECT 11.09 1.22 11.985 1.55 ;
      RECT 11.09 0.54 11.31 1.22 ;
      RECT 0 3.245 12.48 3.415 ;
      RECT 11.54 1.995 11.87 3.245 ;
      RECT 6.45 2.86 6.78 3.245 ;
      RECT 2.56 2.73 3.15 3.245 ;
      RECT 3.83 2.73 4.335 3.245 ;
      RECT 8.86 2.65 9.43 3.245 ;
      RECT 10.12 1.82 10.45 3.245 ;
      RECT 0.7 2.3 1.03 3.245 ;
      RECT 0 -0.085 12.48 0.085 ;
      RECT 11.49 0.085 11.865 1.02 ;
      RECT 2.615 0.085 2.865 0.81 ;
      RECT 3.595 0.085 3.935 0.67 ;
      RECT 6.43 0.085 6.68 0.52 ;
      RECT 8.74 0.085 9.41 0.81 ;
      RECT 10.15 0.085 10.32 1.13 ;
      RECT 0.635 0.085 0.965 0.73 ;
      RECT 5.935 2.52 7.735 2.69 ;
      RECT 5.935 2.2 6.105 2.52 ;
      RECT 7.565 1.96 7.735 2.52 ;
      RECT 5.75 1.87 6.105 2.2 ;
      RECT 7.565 1.63 7.88 1.96 ;
      RECT 0.745 1.955 2.17 2.125 ;
      RECT 1.84 1.795 2.17 1.955 ;
      RECT 0.085 0.785 0.255 1.525 ;
      RECT 0.085 1.855 0.53 2.98 ;
      RECT 0.085 1.525 0.915 1.855 ;
      RECT 0.745 1.855 0.915 1.955 ;
      RECT 0.085 0.35 0.465 0.785 ;
      RECT 4.91 2.22 5.24 2.28 ;
      RECT 4.535 1.82 5.24 2.22 ;
      RECT 5.07 0.425 5.24 1.82 ;
      RECT 4.195 0.255 6.035 0.425 ;
      RECT 4.195 0.425 4.445 1.13 ;
      RECT 5.75 0.425 6.035 0.69 ;
      RECT 5.75 0.69 7.02 0.86 ;
      RECT 5.75 0.86 6.035 1.36 ;
      RECT 6.85 0.425 7.02 0.69 ;
      RECT 6.85 0.255 7.86 0.425 ;
      RECT 7.69 0.425 7.86 1.09 ;
      RECT 7.53 1.09 7.86 1.25 ;
      RECT 7.53 1.25 8.22 1.355 ;
      RECT 7.53 1.355 8.68 1.42 ;
      RECT 8.05 1.42 8.68 1.61 ;
      RECT 3.27 1.99 3.6 2.22 ;
      RECT 3.27 1.82 4.025 1.99 ;
      RECT 3.855 1.01 4.025 1.82 ;
      RECT 3.035 0.84 4.025 1.01 ;
      RECT 3.035 0.35 3.365 0.84 ;
      RECT 7.905 2.13 8.235 2.98 ;
      RECT 8.065 1.95 8.235 2.13 ;
      RECT 8.065 1.78 9.02 1.95 ;
      RECT 8.85 1.27 9.02 1.78 ;
      RECT 8.85 1.15 9.61 1.27 ;
      RECT 9.28 1.27 9.61 1.77 ;
      RECT 8.39 1.1 9.61 1.15 ;
      RECT 8.39 0.98 9.02 1.1 ;
      RECT 8.39 0.81 8.56 0.98 ;
      RECT 8.03 0.35 8.56 0.81 ;
      RECT 4.985 2.63 5.235 2.92 ;
      RECT 4.505 2.56 5.235 2.63 ;
      RECT 1.57 2.46 5.235 2.56 ;
      RECT 1.57 2.39 4.675 2.46 ;
      RECT 4.195 1.65 4.365 2.39 ;
      RECT 4.195 1.48 4.9 1.65 ;
      RECT 4.65 0.595 4.9 1.48 ;
      RECT 2.895 1.35 3.065 2.39 ;
      RECT 2.22 1.18 3.065 1.35 ;
      RECT 2.22 0.64 2.39 1.18 ;
      RECT 1.455 0.39 2.39 0.64 ;
      RECT 1.57 2.56 1.9 2.98 ;
      RECT 1.57 2.3 1.9 2.39 ;
  END
END scs8ls_sdfxbp_1

MACRO scs8ls_sdfxbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.075 1.15 13.315 1.82 ;
        RECT 12.555 1.82 13.315 2.15 ;
        RECT 12.55 0.9 13.315 1.15 ;
        RECT 12.555 2.15 12.835 2.98 ;
    END
    ANTENNADIFFAREA 0.5543 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.62 0.35 10.95 1.13 ;
        RECT 10.78 1.13 10.95 1.8 ;
        RECT 10.59 1.8 10.95 1.97 ;
        RECT 10.59 1.97 10.84 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END Q

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405 1.775 2.755 2.15 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.47 1.655 1.8 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.265 1.35 3.685 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.9 2.075 1.23 ;
        RECT 1.565 0.81 2.075 0.9 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.44 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.44 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
    LAYER li1 ;
      RECT 6.035 2.615 7.735 2.785 ;
      RECT 6.035 2.245 6.205 2.615 ;
      RECT 7.565 1.93 7.735 2.615 ;
      RECT 5.845 1.915 6.205 2.245 ;
      RECT 7.565 1.6 7.895 1.93 ;
      RECT 7.905 2.1 8.235 2.98 ;
      RECT 8.065 1.89 8.235 2.1 ;
      RECT 8.065 1.72 9.02 1.89 ;
      RECT 8.85 1.225 9.02 1.72 ;
      RECT 8.85 1.055 9.61 1.225 ;
      RECT 9.28 1.225 9.61 1.55 ;
      RECT 8.02 0.885 9.02 1.055 ;
      RECT 8.02 0.81 8.19 0.885 ;
      RECT 7.86 0.35 8.19 0.81 ;
      RECT 0.745 1.97 2.195 2.14 ;
      RECT 1.865 1.725 2.195 1.97 ;
      RECT 0.085 0.73 0.255 1.47 ;
      RECT 0.085 1.8 0.52 2.925 ;
      RECT 0.085 1.47 0.915 1.8 ;
      RECT 0.745 1.8 0.915 1.97 ;
      RECT 0.085 0.35 0.49 0.73 ;
      RECT 5.005 2.2 5.335 2.325 ;
      RECT 4.605 2.005 5.335 2.2 ;
      RECT 4.605 1.82 4.855 2.005 ;
      RECT 5.07 0.425 5.24 2.005 ;
      RECT 4.195 0.255 6.08 0.425 ;
      RECT 4.195 0.425 4.445 1.13 ;
      RECT 5.91 0.425 6.08 0.77 ;
      RECT 5.91 0.77 7.01 0.94 ;
      RECT 5.91 0.94 6.08 1.045 ;
      RECT 6.84 0.425 7.01 0.77 ;
      RECT 5.75 1.045 6.08 1.375 ;
      RECT 6.84 0.255 7.69 0.425 ;
      RECT 7.52 0.425 7.69 1.03 ;
      RECT 7.52 1.03 7.78 1.225 ;
      RECT 7.52 1.225 8.68 1.395 ;
      RECT 8.35 1.395 8.68 1.55 ;
      RECT 5.085 2.665 5.335 2.935 ;
      RECT 4.575 2.54 5.335 2.665 ;
      RECT 1.65 2.495 5.335 2.54 ;
      RECT 1.65 2.37 4.745 2.495 ;
      RECT 4.265 1.65 4.435 2.37 ;
      RECT 4.265 1.48 4.9 1.65 ;
      RECT 4.65 0.595 4.9 1.48 ;
      RECT 2.925 1.52 3.095 2.37 ;
      RECT 2.245 1.35 3.095 1.52 ;
      RECT 2.245 0.64 2.415 1.35 ;
      RECT 1.48 0.39 2.415 0.64 ;
      RECT 1.65 2.54 1.98 2.925 ;
      RECT 1.65 2.31 1.98 2.37 ;
      RECT 0 -0.085 13.44 0.085 ;
      RECT 12.995 0.085 13.325 0.73 ;
      RECT 11.13 0.085 11.38 1.13 ;
      RECT 12.12 0.085 12.45 0.73 ;
      RECT 12.12 0.73 12.38 1.15 ;
      RECT 2.695 0.085 2.945 1.13 ;
      RECT 3.685 0.085 4.015 0.84 ;
      RECT 6.34 0.085 6.67 0.6 ;
      RECT 8.68 0.085 9.39 0.715 ;
      RECT 10.12 0.085 10.45 1.13 ;
      RECT 0.66 0.085 0.99 0.73 ;
      RECT 0 3.245 13.44 3.415 ;
      RECT 13.005 2.32 13.335 3.245 ;
      RECT 11.04 2.14 11.37 3.245 ;
      RECT 12.105 1.82 12.355 3.245 ;
      RECT 11.12 1.82 11.37 2.14 ;
      RECT 6.575 2.955 6.905 3.245 ;
      RECT 2.67 2.71 3.09 3.245 ;
      RECT 4.075 2.71 4.405 3.245 ;
      RECT 8.86 2.65 9.43 3.245 ;
      RECT 10.14 1.82 10.39 3.245 ;
      RECT 0.725 2.31 1.055 3.245 ;
      RECT 5.505 2.475 5.865 2.935 ;
      RECT 5.505 1.745 5.675 2.475 ;
      RECT 5.41 1.575 7.01 1.745 ;
      RECT 6.73 1.745 7.01 1.945 ;
      RECT 5.41 0.875 5.58 1.575 ;
      RECT 5.41 0.595 5.74 0.875 ;
      RECT 7.11 2.115 7.395 2.445 ;
      RECT 7.18 1.405 7.35 2.115 ;
      RECT 6.25 1.11 7.35 1.405 ;
      RECT 7.18 0.595 7.35 1.11 ;
      RECT 3.295 1.95 4.095 2.2 ;
      RECT 3.855 1.35 4.095 1.95 ;
      RECT 3.855 1.18 4.025 1.35 ;
      RECT 3.125 1.01 4.025 1.18 ;
      RECT 3.125 0.35 3.455 1.01 ;
      RECT 11.58 1.32 12.735 1.65 ;
      RECT 11.58 1.65 11.91 2.86 ;
      RECT 11.58 0.56 11.94 1.32 ;
      RECT 9.78 1.3 10.61 1.63 ;
      RECT 9.6 2.38 9.95 2.98 ;
      RECT 8.71 2.06 9.95 2.38 ;
      RECT 9.6 1.94 9.95 2.06 ;
      RECT 9.78 1.63 9.95 1.94 ;
      RECT 9.78 0.885 9.95 1.3 ;
      RECT 9.56 0.35 9.95 0.885 ;
  END
END scs8ls_sdfxbp_2

MACRO scs8ls_sdfxtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 11.04 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.455 1.655 1.785 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405 1.47 2.74 2.14 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.25 1.18 3.685 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.6 0.37 10.935 2.98 ;
    END
    ANTENNADIFFAREA 0.5283 ;
  END Q

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 0.9 2.25 0.955 ;
        RECT 0.425 0.955 2.25 1.285 ;
        RECT 1.085 0.81 1.315 0.9 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.04 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.04 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
    LAYER li1 ;
      RECT 0 -0.085 11.04 0.085 ;
      RECT 2.775 0.085 2.945 0.79 ;
      RECT 3.685 0.085 4.015 0.62 ;
      RECT 6.385 0.085 6.635 0.52 ;
      RECT 8.805 0.085 9.48 0.81 ;
      RECT 10.175 0.085 10.425 1.15 ;
      RECT 0.585 0.085 0.915 0.785 ;
      RECT 7.015 2.1 7.375 2.35 ;
      RECT 7.145 1.36 7.315 2.1 ;
      RECT 6.195 1.03 7.315 1.36 ;
      RECT 7.145 0.86 7.315 1.03 ;
      RECT 7.145 0.595 7.475 0.86 ;
      RECT 4.955 2.22 5.225 2.38 ;
      RECT 4.565 2.05 5.225 2.22 ;
      RECT 4.565 1.82 4.815 2.05 ;
      RECT 5.055 0.425 5.225 2.05 ;
      RECT 4.195 0.255 5.905 0.425 ;
      RECT 4.195 0.425 4.445 1.13 ;
      RECT 5.735 0.425 5.905 0.69 ;
      RECT 5.735 0.69 6.975 0.86 ;
      RECT 5.735 0.86 5.985 1.36 ;
      RECT 6.805 0.425 6.975 0.69 ;
      RECT 6.805 0.255 7.815 0.425 ;
      RECT 7.645 0.425 7.815 1.03 ;
      RECT 7.485 1.03 7.815 1.19 ;
      RECT 7.485 1.19 8.24 1.32 ;
      RECT 7.485 1.32 8.555 1.36 ;
      RECT 8.07 1.36 8.555 1.49 ;
      RECT 8.305 1.49 8.555 2.075 ;
      RECT 6.045 2.52 7.715 2.69 ;
      RECT 6.045 2.2 6.215 2.52 ;
      RECT 7.545 1.93 7.715 2.52 ;
      RECT 5.735 1.87 6.215 2.2 ;
      RECT 7.545 1.6 7.9 1.93 ;
      RECT 3.295 1.82 4.055 2.14 ;
      RECT 3.855 1.3 4.055 1.82 ;
      RECT 3.855 0.96 4.025 1.3 ;
      RECT 3.125 0.79 4.025 0.96 ;
      RECT 3.125 0.35 3.455 0.79 ;
      RECT 7.885 2.415 8.135 2.98 ;
      RECT 7.885 2.245 8.895 2.415 ;
      RECT 7.885 2.1 8.135 2.245 ;
      RECT 8.725 1.93 8.895 2.245 ;
      RECT 8.725 1.6 9.595 1.93 ;
      RECT 8.725 1.15 8.895 1.6 ;
      RECT 8.41 0.98 8.895 1.15 ;
      RECT 8.41 0.94 8.58 0.98 ;
      RECT 7.985 0.77 8.58 0.94 ;
      RECT 7.985 0.48 8.315 0.77 ;
      RECT 0.085 1.955 2.195 2.125 ;
      RECT 1.865 2.125 2.195 2.14 ;
      RECT 1.865 1.47 2.195 1.955 ;
      RECT 0.085 0.785 0.255 1.525 ;
      RECT 0.085 0.35 0.405 0.785 ;
      RECT 0.085 2.125 0.555 2.98 ;
      RECT 0.085 1.525 0.825 1.955 ;
      RECT 4.535 2.71 5.375 2.98 ;
      RECT 4.535 2.56 4.705 2.71 ;
      RECT 3.345 2.48 4.705 2.56 ;
      RECT 1.595 2.39 4.705 2.48 ;
      RECT 1.595 2.31 4.395 2.39 ;
      RECT 4.225 1.65 4.395 2.31 ;
      RECT 4.225 1.48 4.785 1.65 ;
      RECT 4.615 0.94 4.785 1.48 ;
      RECT 4.615 0.595 4.885 0.94 ;
      RECT 2.91 1.3 3.08 2.31 ;
      RECT 2.42 1.13 3.08 1.3 ;
      RECT 2.42 0.73 2.59 1.13 ;
      RECT 1.485 0.4 2.59 0.73 ;
      RECT 1.595 2.48 1.925 2.98 ;
      RECT 5.545 2.54 5.875 2.98 ;
      RECT 5.395 2.37 5.875 2.54 ;
      RECT 5.395 1.7 5.565 2.37 ;
      RECT 5.395 1.53 6.975 1.7 ;
      RECT 6.645 1.7 6.975 1.93 ;
      RECT 5.395 0.595 5.565 1.53 ;
      RECT 9.59 2.1 9.935 2.98 ;
      RECT 9.765 1.65 9.935 2.1 ;
      RECT 9.765 1.36 10.245 1.65 ;
      RECT 9.065 1.32 10.245 1.36 ;
      RECT 9.065 1.03 9.98 1.32 ;
      RECT 9.65 0.35 9.98 1.03 ;
      RECT 0 3.245 11.04 3.415 ;
      RECT 6.48 2.86 6.81 3.245 ;
      RECT 3.855 2.73 4.365 3.245 ;
      RECT 2.67 2.65 3.175 3.245 ;
      RECT 8.845 2.65 9.42 3.245 ;
      RECT 10.15 1.82 10.4 3.245 ;
      RECT 0.725 2.3 1.055 3.245 ;
  END
END scs8ls_sdfxtp_1

MACRO scs8ls_sdfxtp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.105 1.82 11.435 2.98 ;
        RECT 11.215 1.05 11.385 1.82 ;
        RECT 11.055 0.35 11.385 1.05 ;
    END
    ANTENNADIFFAREA 0.5765 ;
  END Q

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.45 1.435 2.78 2.15 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.19 1.665 1.845 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.29 1.35 3.685 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.85 2.205 1.02 ;
        RECT 0.425 1.02 0.835 1.23 ;
        RECT 1.875 1.02 2.205 1.23 ;
        RECT 0.425 0.81 0.835 0.85 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
    LAYER li1 ;
      RECT 0 3.245 12 3.415 ;
      RECT 11.635 1.82 11.885 3.245 ;
      RECT 2.685 2.79 3.135 3.245 ;
      RECT 3.9 2.79 4.37 3.245 ;
      RECT 9.295 2.59 9.925 3.245 ;
      RECT 6.585 2.52 6.835 3.245 ;
      RECT 10.655 1.82 10.905 3.245 ;
      RECT 0.615 2.355 0.945 3.245 ;
      RECT 7.005 2.905 7.855 3.075 ;
      RECT 7.005 2.3 7.175 2.905 ;
      RECT 7.685 1.93 7.855 2.905 ;
      RECT 5.895 2.13 7.175 2.3 ;
      RECT 7.685 1.6 8.115 1.93 ;
      RECT 5.895 1.97 6.225 2.13 ;
      RECT 7.345 1.39 7.515 2.61 ;
      RECT 6.485 1.23 7.515 1.39 ;
      RECT 6.485 1.06 7.89 1.23 ;
      RECT 7.56 0.595 7.89 1.06 ;
      RECT 8.285 1.99 8.72 2.32 ;
      RECT 8.285 1.36 8.455 1.99 ;
      RECT 8.06 1.03 8.455 1.36 ;
      RECT 8.06 0.425 8.23 1.03 ;
      RECT 7.22 0.255 8.23 0.425 ;
      RECT 7.22 0.425 7.39 0.72 ;
      RECT 5.945 0.72 7.39 0.89 ;
      RECT 5.945 0.89 6.275 1.36 ;
      RECT 5.945 0.425 6.115 0.72 ;
      RECT 4.205 0.255 6.115 0.425 ;
      RECT 4.205 0.425 4.535 1.13 ;
      RECT 5.185 0.425 5.355 1.61 ;
      RECT 5.045 1.61 5.375 1.82 ;
      RECT 4.655 1.82 5.375 2.28 ;
      RECT 8.025 2.66 8.275 2.92 ;
      RECT 8.025 2.49 9.06 2.66 ;
      RECT 8.89 2.245 9.06 2.49 ;
      RECT 8.89 2.075 10.105 2.245 ;
      RECT 9.775 1.41 10.105 2.075 ;
      RECT 8.89 0.81 9.06 2.075 ;
      RECT 8.4 0.64 9.06 0.81 ;
      RECT 8.4 0.35 8.795 0.64 ;
      RECT 0.085 2.015 2.21 2.185 ;
      RECT 1.88 1.775 2.21 2.015 ;
      RECT 0.085 0.64 0.255 1.47 ;
      RECT 0.085 2.185 0.445 2.925 ;
      RECT 0.085 1.47 0.915 2.015 ;
      RECT 0.085 0.39 0.49 0.64 ;
      RECT 1.485 2.45 5.385 2.62 ;
      RECT 5.135 2.62 5.385 2.98 ;
      RECT 4.315 1.47 4.485 2.45 ;
      RECT 4.315 1.3 4.875 1.47 ;
      RECT 4.705 0.94 4.875 1.3 ;
      RECT 4.705 0.595 5.015 0.94 ;
      RECT 1.485 2.355 3.12 2.45 ;
      RECT 2.95 1.265 3.12 2.355 ;
      RECT 2.375 1.095 3.12 1.265 ;
      RECT 2.375 0.68 2.545 1.095 ;
      RECT 1.48 0.35 2.545 0.68 ;
      RECT 1.485 2.62 2.06 2.945 ;
      RECT 3.34 1.95 4.145 2.28 ;
      RECT 3.855 1.3 4.145 1.95 ;
      RECT 3.855 1.18 4.025 1.3 ;
      RECT 3.305 1.01 4.025 1.18 ;
      RECT 3.305 0.92 3.475 1.01 ;
      RECT 3.145 0.33 3.475 0.92 ;
      RECT 5.555 2.52 5.915 2.98 ;
      RECT 5.555 1.8 5.725 2.52 ;
      RECT 5.555 1.63 7.175 1.8 ;
      RECT 6.845 1.8 7.175 1.96 ;
      RECT 5.555 0.94 5.775 1.63 ;
      RECT 5.525 0.595 5.775 0.94 ;
      RECT 10.095 2.415 10.445 2.92 ;
      RECT 10.275 1.55 10.445 2.415 ;
      RECT 10.275 1.24 11.045 1.55 ;
      RECT 9.23 1.22 11.045 1.24 ;
      RECT 9.23 1.24 9.535 1.905 ;
      RECT 9.23 1.07 10.445 1.22 ;
      RECT 9.8 0.35 10.13 1.07 ;
      RECT 0 -0.085 12 0.085 ;
      RECT 11.555 0.085 11.885 1.13 ;
      RECT 2.715 0.085 2.975 0.81 ;
      RECT 3.705 0.085 4.035 0.84 ;
      RECT 6.72 0.085 7.05 0.55 ;
      RECT 9.3 0.085 9.63 0.81 ;
      RECT 10.615 0.085 10.885 1.05 ;
      RECT 0.66 0.085 0.99 0.64 ;
  END
END scs8ls_sdfxtp_2

MACRO scs8ls_sdfxtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.48 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.76 1.13 12.355 1.8 ;
        RECT 10.685 1.8 12.355 1.97 ;
        RECT 10.745 0.88 12.355 1.13 ;
        RECT 11.665 1.97 12.355 2.015 ;
        RECT 10.685 1.97 11.015 2.98 ;
        RECT 10.745 0.35 10.995 0.88 ;
        RECT 11.675 0.35 11.865 0.88 ;
        RECT 11.665 2.015 11.855 2.98 ;
    END
    ANTENNADIFFAREA 1.1493 ;
  END Q

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.435 1.55 2.765 2.15 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.455 1.655 1.785 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.275 1.18 3.685 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.81 2.195 0.955 ;
        RECT 0.425 0.955 2.195 1.285 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12.48 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12.48 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
    LAYER li1 ;
      RECT 0 -0.085 12.48 0.085 ;
      RECT 12.035 0.085 12.365 0.71 ;
      RECT 2.705 0.085 2.955 0.81 ;
      RECT 3.685 0.085 4.015 0.67 ;
      RECT 6.49 0.085 6.82 0.6 ;
      RECT 9.195 0.085 9.525 0.73 ;
      RECT 10.185 0.085 10.515 0.96 ;
      RECT 11.175 0.085 11.505 0.71 ;
      RECT 0.66 0.085 0.99 0.785 ;
      RECT 0 3.245 12.48 3.415 ;
      RECT 12.035 2.185 12.365 3.245 ;
      RECT 6.68 2.855 7.01 3.245 ;
      RECT 2.585 2.73 3.205 3.245 ;
      RECT 3.885 2.73 4.475 3.245 ;
      RECT 9.225 2.36 9.555 3.245 ;
      RECT 10.305 1.94 10.475 3.245 ;
      RECT 11.215 2.14 11.465 3.245 ;
      RECT 0.725 2.3 1.055 3.245 ;
      RECT 9.965 1.3 11.545 1.63 ;
      RECT 9.73 1.97 10.135 2.82 ;
      RECT 9.965 1.63 10.135 1.97 ;
      RECT 9.355 1.13 10.135 1.3 ;
      RECT 9.355 0.9 9.665 1.13 ;
      RECT 9.835 0.35 10.005 1.13 ;
      RECT 6.105 2.515 8.1 2.685 ;
      RECT 6.105 2.28 6.275 2.515 ;
      RECT 7.93 1.955 8.1 2.515 ;
      RECT 5.915 1.95 6.275 2.28 ;
      RECT 7.77 1.625 8.1 1.955 ;
      RECT 7.215 2.175 7.76 2.345 ;
      RECT 7.33 1.44 7.5 2.175 ;
      RECT 6.295 1.11 7.5 1.44 ;
      RECT 7.33 0.885 7.5 1.11 ;
      RECT 7.33 0.635 7.785 0.885 ;
      RECT 5.575 2.51 5.935 2.97 ;
      RECT 5.575 1.78 5.745 2.51 ;
      RECT 5.435 1.61 7.16 1.78 ;
      RECT 6.835 1.78 7.16 1.94 ;
      RECT 5.435 0.595 5.605 1.61 ;
      RECT 5.155 2.71 5.405 2.97 ;
      RECT 4.645 2.56 5.405 2.71 ;
      RECT 1.595 2.54 5.405 2.56 ;
      RECT 1.595 2.39 4.815 2.54 ;
      RECT 4.335 1.65 4.505 2.39 ;
      RECT 4.335 1.48 4.925 1.65 ;
      RECT 4.675 0.595 4.925 1.48 ;
      RECT 2.935 1.35 3.105 2.39 ;
      RECT 2.365 1.18 3.105 1.35 ;
      RECT 2.365 0.64 2.535 1.18 ;
      RECT 1.48 0.39 2.535 0.64 ;
      RECT 1.595 2.56 1.925 2.98 ;
      RECT 1.595 2.31 1.925 2.39 ;
      RECT 8.27 2.19 8.6 2.82 ;
      RECT 8.27 2.02 9.185 2.19 ;
      RECT 9.015 1.8 9.185 2.02 ;
      RECT 9.015 1.47 9.795 1.8 ;
      RECT 9.015 1.07 9.185 1.47 ;
      RECT 8.295 0.9 9.185 1.07 ;
      RECT 8.295 0.35 8.625 0.9 ;
      RECT 0.085 1.955 2.195 2.125 ;
      RECT 1.865 2.125 2.195 2.14 ;
      RECT 1.865 1.47 2.195 1.955 ;
      RECT 0.085 0.785 0.255 1.525 ;
      RECT 0.085 2.125 0.555 2.98 ;
      RECT 0.085 1.525 0.915 1.955 ;
      RECT 0.085 0.35 0.49 0.785 ;
      RECT 3.325 1.99 3.655 2.22 ;
      RECT 3.325 1.82 4.165 1.99 ;
      RECT 3.855 1.3 4.165 1.82 ;
      RECT 3.855 1.01 4.025 1.3 ;
      RECT 3.125 0.84 4.025 1.01 ;
      RECT 3.125 0.35 3.455 0.84 ;
      RECT 5.075 2.22 5.405 2.37 ;
      RECT 4.675 2.04 5.405 2.22 ;
      RECT 4.675 1.82 4.925 2.04 ;
      RECT 5.095 0.425 5.265 2.04 ;
      RECT 4.195 0.255 5.945 0.425 ;
      RECT 4.195 0.425 4.445 1.13 ;
      RECT 5.775 0.425 5.945 0.77 ;
      RECT 5.775 0.77 7.16 0.94 ;
      RECT 5.775 0.94 6.075 1.36 ;
      RECT 6.99 0.465 7.16 0.77 ;
      RECT 6.99 0.295 8.125 0.465 ;
      RECT 7.955 0.465 8.125 1.055 ;
      RECT 7.67 1.055 8.125 1.24 ;
      RECT 7.67 1.24 8.845 1.41 ;
      RECT 8.535 1.41 8.845 1.715 ;
  END
END scs8ls_sdfxtp_4

MACRO scs8ls_sdlclkp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.29 0.545 1.96 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END SCE

  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805 1.63 1.285 2.15 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END GATE

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 5.33 1.355 5.66 1.78 ;
    END
    ANTENNAGATEAREA 0.459 ;
  END CLK

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.235 1.82 7.585 2.98 ;
        RECT 7.415 1.13 7.585 1.82 ;
        RECT 7.24 0.35 7.585 1.13 ;
    END
    ANTENNADIFFAREA 0.6328 ;
  END GCLK

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.795 1.715 2.38 2.15 ;
      RECT 1.795 1.545 2.9 1.715 ;
      RECT 2.625 1.385 2.9 1.545 ;
      RECT 1.795 1.12 1.965 1.545 ;
      RECT 1.565 0.95 1.965 1.12 ;
      RECT 1.565 0.88 1.895 0.95 ;
      RECT 6.475 1.3 7.245 1.63 ;
      RECT 6.195 1.89 6.525 2.875 ;
      RECT 6.195 1.72 6.645 1.89 ;
      RECT 6.475 1.63 6.645 1.72 ;
      RECT 6.475 1.05 6.645 1.3 ;
      RECT 6.165 0.45 6.645 1.05 ;
      RECT 4.49 2.495 6 2.665 ;
      RECT 5.83 1.55 6 2.495 ;
      RECT 5.83 1.22 6.305 1.55 ;
      RECT 4.49 2.665 4.82 2.9 ;
      RECT 4.49 2.12 4.82 2.495 ;
      RECT 3.6 1.74 4.82 2.12 ;
      RECT 4.49 1.05 4.68 1.74 ;
      RECT 4.43 0.595 4.68 1.05 ;
      RECT 4.99 1.995 5.38 2.325 ;
      RECT 4.99 1.13 5.16 1.995 ;
      RECT 4.9 0.425 5.23 1.13 ;
      RECT 4.09 0.255 5.23 0.425 ;
      RECT 4.09 0.425 4.26 0.88 ;
      RECT 3.41 0.88 4.26 1.05 ;
      RECT 3.41 0.425 3.58 0.88 ;
      RECT 2.545 0.255 3.58 0.425 ;
      RECT 2.545 0.425 2.715 1.03 ;
      RECT 2.135 1.03 2.715 1.2 ;
      RECT 2.135 1.2 2.415 1.36 ;
      RECT 3.06 2.425 3.39 2.755 ;
      RECT 3.07 1.55 3.39 2.425 ;
      RECT 3.07 1.22 4.32 1.55 ;
      RECT 3.07 0.925 3.24 1.22 ;
      RECT 2.885 0.595 3.24 0.925 ;
      RECT 0.955 2.49 1.285 2.98 ;
      RECT 0.955 2.32 2.86 2.49 ;
      RECT 2.61 2.49 2.86 2.755 ;
      RECT 2.61 1.885 2.86 2.32 ;
      RECT 1.455 1.46 1.625 2.32 ;
      RECT 0.715 1.29 1.625 1.46 ;
      RECT 0.715 1.12 0.885 1.29 ;
      RECT 0.545 0.71 0.885 1.12 ;
      RECT 0.545 0.54 2.375 0.71 ;
      RECT 2.125 0.71 2.375 0.78 ;
      RECT 2.125 0.35 2.375 0.54 ;
      RECT 0 3.245 7.68 3.415 ;
      RECT 5.585 2.835 5.99 3.245 ;
      RECT 1.515 2.66 1.845 3.245 ;
      RECT 3.985 2.44 4.315 3.245 ;
      RECT 6.695 2.06 7.025 3.245 ;
      RECT 0.115 2.13 0.445 3.245 ;
      RECT 0 -0.085 7.68 0.085 ;
      RECT 0.115 0.085 0.365 1.12 ;
      RECT 1.055 0.085 1.385 0.37 ;
      RECT 3.75 0.085 3.92 0.71 ;
      RECT 5.41 0.085 5.66 1.13 ;
      RECT 6.815 0.085 7.065 1.13 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
  END
END scs8ls_sdlclkp_1

MACRO scs8ls_sdlclkp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.29 0.55 1.96 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END SCE

  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.795 1.63 1.3 2.15 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END GATE

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 5.335 1.18 5.665 1.55 ;
    END
    ANTENNAGATEAREA 0.498 ;
  END CLK

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.21 1.82 7.565 2.98 ;
        RECT 7.395 1.13 7.565 1.82 ;
        RECT 7.295 0.35 7.625 1.13 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END GCLK

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.81 1.715 2.34 2.15 ;
      RECT 1.81 1.545 3.02 1.715 ;
      RECT 2.69 1.385 3.02 1.545 ;
      RECT 1.81 1.05 1.98 1.545 ;
      RECT 1.565 0.88 1.98 1.05 ;
      RECT 4.44 2.22 6.005 2.39 ;
      RECT 5.835 1.63 6.005 2.22 ;
      RECT 5.835 1.3 6.53 1.63 ;
      RECT 4.44 2.39 4.825 2.92 ;
      RECT 4.44 1.925 4.825 2.22 ;
      RECT 3.53 1.755 4.825 1.925 ;
      RECT 3.53 1.585 3.86 1.755 ;
      RECT 4.655 1.075 4.825 1.755 ;
      RECT 4.55 0.595 4.825 1.075 ;
      RECT 3 2.235 3.36 2.695 ;
      RECT 3.19 1.415 3.36 2.235 ;
      RECT 3.19 1.245 4.485 1.415 ;
      RECT 4.155 1.415 4.485 1.585 ;
      RECT 3.19 0.845 3.36 1.245 ;
      RECT 2.885 0.595 3.36 0.845 ;
      RECT 0.945 2.49 1.275 2.98 ;
      RECT 0.945 2.32 2.8 2.49 ;
      RECT 2.55 2.49 2.8 2.755 ;
      RECT 2.55 1.885 2.8 2.32 ;
      RECT 1.47 1.39 1.64 2.32 ;
      RECT 0.72 1.22 1.64 1.39 ;
      RECT 0.72 1.12 0.89 1.22 ;
      RECT 0.545 0.71 0.89 1.12 ;
      RECT 0.545 0.54 2.375 0.71 ;
      RECT 2.125 0.35 2.375 0.54 ;
      RECT 4.995 0.425 5.36 1.01 ;
      RECT 4.21 0.255 5.36 0.425 ;
      RECT 4.995 1.72 5.31 2.05 ;
      RECT 4.995 1.01 5.165 1.72 ;
      RECT 4.21 0.425 4.38 0.905 ;
      RECT 3.53 0.905 4.38 1.075 ;
      RECT 3.53 0.425 3.7 0.905 ;
      RECT 2.545 0.255 3.7 0.425 ;
      RECT 2.545 0.425 2.715 1.03 ;
      RECT 2.15 1.03 2.715 1.2 ;
      RECT 2.15 1.2 2.48 1.36 ;
      RECT 6.87 1.3 7.225 1.63 ;
      RECT 6.175 1.97 6.505 2.89 ;
      RECT 6.175 1.8 7.04 1.97 ;
      RECT 6.87 1.63 7.04 1.8 ;
      RECT 6.87 1.13 7.04 1.3 ;
      RECT 6.325 0.96 7.04 1.13 ;
      RECT 6.325 0.35 6.655 0.96 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 7.74 1.82 7.99 3.245 ;
      RECT 1.485 2.66 1.815 3.245 ;
      RECT 5.51 2.56 5.84 3.245 ;
      RECT 6.71 2.14 7.04 3.245 ;
      RECT 3.99 2.095 4.24 3.245 ;
      RECT 0.105 2.13 0.435 3.245 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 7.805 0.085 8.055 1.13 ;
      RECT 0.115 0.085 0.365 1.12 ;
      RECT 1.055 0.085 1.385 0.37 ;
      RECT 3.87 0.085 4.04 0.735 ;
      RECT 5.53 0.085 5.86 1.01 ;
      RECT 6.865 0.085 7.115 0.79 ;
    LAYER mcon ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
  END
END scs8ls_sdlclkp_2

MACRO scs8ls_sdlclkp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.725 1.13 9.055 1.41 ;
        RECT 8.725 1.41 8.985 1.8 ;
        RECT 7.865 0.96 9.055 1.13 ;
        RECT 7.705 1.8 8.985 1.97 ;
        RECT 7.865 0.35 8.115 0.96 ;
        RECT 8.725 0.35 9.055 0.96 ;
        RECT 7.705 1.97 8.035 2.98 ;
        RECT 8.655 1.97 8.985 2.98 ;
    END
    ANTENNADIFFAREA 1.3194 ;
  END GCLK

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 5.785 1.18 6.115 1.55 ;
    END
    ANTENNAGATEAREA 0.516 ;
  END CLK

  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835 1.455 1.315 1.785 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END GATE

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.455 0.55 1.785 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END SCE

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.365 1.735 2.695 2.14 ;
      RECT 1.825 1.565 3.255 1.735 ;
      RECT 2.925 1.405 3.255 1.565 ;
      RECT 1.825 0.955 2.075 1.565 ;
      RECT 0.985 2.48 1.315 2.835 ;
      RECT 0.985 2.31 3.255 2.48 ;
      RECT 2.925 2.48 3.255 2.755 ;
      RECT 0.985 1.955 1.655 2.31 ;
      RECT 2.925 1.905 3.255 2.31 ;
      RECT 1.485 0.785 1.655 1.955 ;
      RECT 0.615 0.615 2.635 0.785 ;
      RECT 0.615 0.785 0.945 1.285 ;
      RECT 2.305 0.785 2.635 0.895 ;
      RECT 2.305 0.35 2.635 0.615 ;
      RECT 5.445 0.425 5.835 1.01 ;
      RECT 4.605 0.255 5.835 0.425 ;
      RECT 5.44 1.82 5.775 2.07 ;
      RECT 5.445 1.01 5.615 1.82 ;
      RECT 4.605 0.425 4.775 0.895 ;
      RECT 3.765 0.895 4.775 1.065 ;
      RECT 3.765 0.44 3.935 0.895 ;
      RECT 2.805 0.27 3.935 0.44 ;
      RECT 2.805 0.44 2.975 1.065 ;
      RECT 2.245 1.065 2.975 1.235 ;
      RECT 2.245 1.235 2.575 1.395 ;
      RECT 4.88 2.24 6.455 2.41 ;
      RECT 6.285 1.63 6.455 2.24 ;
      RECT 6.285 1.3 7.03 1.63 ;
      RECT 4.88 2.41 5.27 2.895 ;
      RECT 4.88 1.905 5.27 2.24 ;
      RECT 3.96 1.735 5.27 1.905 ;
      RECT 3.96 1.575 4.29 1.735 ;
      RECT 5.1 1.065 5.27 1.735 ;
      RECT 4.945 0.595 5.275 1.065 ;
      RECT 3.425 1.405 3.705 2.755 ;
      RECT 3.425 1.235 4.93 1.405 ;
      RECT 4.6 1.405 4.93 1.565 ;
      RECT 3.425 0.94 3.595 1.235 ;
      RECT 3.145 0.61 3.595 0.94 ;
      RECT 7.365 1.3 8.435 1.63 ;
      RECT 6.625 1.97 6.955 2.98 ;
      RECT 6.625 1.8 7.535 1.97 ;
      RECT 7.365 1.63 7.535 1.8 ;
      RECT 7.365 1.13 7.535 1.3 ;
      RECT 6.825 0.96 7.535 1.13 ;
      RECT 6.825 0.35 7.155 0.96 ;
      RECT 0 3.245 9.6 3.415 ;
      RECT 9.155 1.82 9.485 3.245 ;
      RECT 1.545 2.65 2.16 3.245 ;
      RECT 5.98 2.58 6.31 3.245 ;
      RECT 7.125 2.14 7.455 3.245 ;
      RECT 4.43 2.075 4.68 3.245 ;
      RECT 0.115 1.955 0.445 3.245 ;
      RECT 8.235 2.14 8.485 3.245 ;
      RECT 0 -0.085 9.6 0.085 ;
      RECT 9.235 0.085 9.485 1.13 ;
      RECT 6.005 0.085 6.335 1.01 ;
      RECT 7.385 0.085 7.635 0.79 ;
      RECT 8.295 0.085 8.545 0.79 ;
      RECT 0.115 0.085 0.445 1.285 ;
      RECT 1.125 0.085 1.565 0.445 ;
      RECT 4.105 0.085 4.435 0.725 ;
    LAYER mcon ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
  END
END scs8ls_sdlclkp_4

MACRO scs8ls_sedfxbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 16.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455 1.06 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.45 2.085 1.78 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END DE

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.475 1.45 4.865 1.78 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.075 1.18 5.635 1.51 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.845 1.82 15.24 2.98 ;
        RECT 14.845 0.62 15.015 1.82 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.575 1.18 7.075 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.86 1.82 16.235 2.98 ;
        RECT 16.065 1.15 16.235 1.82 ;
        RECT 15.875 0.37 16.235 1.15 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END QN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 16.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 16.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 14.075 1.95 14.245 2.12 ;
      RECT 3.035 1.95 3.205 2.12 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
    LAYER met1 ;
      RECT 2.975 2.105 3.265 2.15 ;
      RECT 2.975 1.965 14.305 2.105 ;
      RECT 14.015 2.105 14.305 2.15 ;
      RECT 2.975 1.92 3.265 1.965 ;
      RECT 14.015 1.92 14.305 1.965 ;
    LAYER li1 ;
      RECT 9.19 2.56 9.52 2.98 ;
      RECT 9.04 2.39 9.52 2.56 ;
      RECT 9.04 1.79 9.21 2.39 ;
      RECT 9.04 1.62 10.73 1.79 ;
      RECT 10.4 1.79 10.73 1.83 ;
      RECT 10.4 1.53 10.73 1.62 ;
      RECT 9.04 0.95 9.21 1.62 ;
      RECT 9.04 0.62 9.32 0.95 ;
      RECT 10.615 2.05 11.07 2.22 ;
      RECT 10.9 1.52 11.07 2.05 ;
      RECT 10.9 1.36 11.74 1.52 ;
      RECT 9.86 1.19 11.74 1.36 ;
      RECT 9.86 1.36 10.19 1.45 ;
      RECT 10.9 0.595 11.07 1.19 ;
      RECT 4.055 1.95 5.87 2.12 ;
      RECT 5.565 1.79 5.87 1.95 ;
      RECT 4.055 0.605 4.74 1.065 ;
      RECT 4.135 2.29 4.445 2.735 ;
      RECT 4.135 2.12 4.305 2.29 ;
      RECT 4.055 1.065 4.305 1.95 ;
      RECT 4.055 0.41 4.305 0.605 ;
      RECT 9.69 2.39 12.595 2.56 ;
      RECT 9.69 2.22 9.86 2.39 ;
      RECT 12.425 1.8 12.595 2.39 ;
      RECT 9.38 1.96 9.86 2.22 ;
      RECT 12.425 1.47 12.855 1.8 ;
      RECT 12.765 2.52 13.195 2.98 ;
      RECT 13.025 1.885 13.195 2.52 ;
      RECT 13.025 1.715 13.875 1.885 ;
      RECT 13.705 1.53 13.875 1.715 ;
      RECT 13.705 1.2 14.26 1.53 ;
      RECT 13.705 0.94 13.875 1.2 ;
      RECT 12.29 0.77 13.875 0.94 ;
      RECT 12.29 0.35 12.62 0.77 ;
      RECT 15.185 1.32 15.895 1.65 ;
      RECT 14.205 0.255 15.355 0.425 ;
      RECT 15.185 0.425 15.355 1.32 ;
      RECT 14.43 2.38 14.6 2.98 ;
      RECT 13.46 2.055 14.6 2.38 ;
      RECT 14.045 1.92 14.6 2.055 ;
      RECT 14.43 1.03 14.6 1.92 ;
      RECT 14.205 0.425 14.6 1.03 ;
      RECT 1.375 2.905 2.225 3.075 ;
      RECT 2.055 2.48 2.225 2.905 ;
      RECT 2.055 2.31 3.545 2.48 ;
      RECT 3.185 2.48 3.545 2.98 ;
      RECT 3.375 1.345 3.545 2.31 ;
      RECT 3.03 1.175 3.545 1.345 ;
      RECT 3.03 0.545 3.36 1.175 ;
      RECT 1.375 2.46 1.545 2.905 ;
      RECT 0.115 2.29 1.545 2.46 ;
      RECT 0.115 0.48 0.66 0.81 ;
      RECT 0.115 2.46 0.445 2.98 ;
      RECT 0.115 0.81 0.285 2.29 ;
      RECT 6.725 1.82 7.525 2.14 ;
      RECT 7.055 1.81 7.525 1.82 ;
      RECT 7.355 1.01 7.525 1.81 ;
      RECT 6.73 0.84 7.525 1.01 ;
      RECT 6.73 0.35 7.06 0.84 ;
      RECT 2.875 1.525 3.205 2.14 ;
      RECT 1.715 2.12 1.885 2.735 ;
      RECT 1.025 1.95 2.665 2.12 ;
      RECT 2.335 1.525 2.665 1.95 ;
      RECT 1.025 1.11 2.04 1.28 ;
      RECT 1.71 0.545 2.04 1.11 ;
      RECT 1.025 1.28 1.355 1.95 ;
      RECT 4.615 2.31 8.335 2.46 ;
      RECT 5.715 2.46 8.335 2.48 ;
      RECT 7.775 1.65 7.945 2.31 ;
      RECT 8.165 2.48 8.335 2.73 ;
      RECT 7.775 1.48 8.53 1.65 ;
      RECT 8.165 2.73 9.02 2.98 ;
      RECT 8.28 0.595 8.53 1.48 ;
      RECT 4.615 2.29 6.21 2.31 ;
      RECT 5.715 2.48 6.045 2.97 ;
      RECT 6.04 1.01 6.21 2.29 ;
      RECT 5.74 0.605 6.21 1.01 ;
      RECT 3.715 2.905 4.785 3.075 ;
      RECT 4.615 2.46 4.785 2.905 ;
      RECT 3.715 2.3 3.965 2.905 ;
      RECT 3.715 1.005 3.885 2.3 ;
      RECT 3.53 0.545 3.885 1.005 ;
      RECT 8.585 2.14 8.87 2.38 ;
      RECT 8.115 1.82 8.87 2.14 ;
      RECT 8.7 0.425 8.87 1.82 ;
      RECT 7.8 0.255 9.69 0.425 ;
      RECT 7.8 0.425 8.05 1.13 ;
      RECT 9.49 0.425 9.69 0.85 ;
      RECT 9.49 0.85 10.73 1.02 ;
      RECT 9.49 1.02 9.69 1.12 ;
      RECT 10.56 0.425 10.73 0.85 ;
      RECT 9.38 1.12 9.69 1.45 ;
      RECT 10.56 0.255 11.41 0.425 ;
      RECT 11.24 0.425 11.41 0.85 ;
      RECT 11.24 0.85 12.12 1.02 ;
      RECT 11.95 1.02 12.12 1.13 ;
      RECT 11.95 1.13 13.395 1.3 ;
      RECT 11.95 1.3 12.255 1.8 ;
      RECT 13.065 1.3 13.395 1.545 ;
      RECT 0 -0.085 16.32 0.085 ;
      RECT 15.525 0.085 15.695 1.15 ;
      RECT 1.15 0.085 1.48 0.89 ;
      RECT 2.21 0.085 2.54 1.005 ;
      RECT 4.91 0.085 5.24 1.01 ;
      RECT 6.38 0.085 6.55 1.01 ;
      RECT 7.29 0.085 7.62 0.67 ;
      RECT 10.065 0.085 10.39 0.68 ;
      RECT 11.58 0.085 11.83 0.68 ;
      RECT 13.19 0.085 14.035 0.6 ;
      RECT 0 3.245 16.32 3.415 ;
      RECT 15.44 1.82 15.69 3.245 ;
      RECT 10.08 2.73 10.41 3.245 ;
      RECT 11.175 2.73 11.505 3.245 ;
      RECT 2.395 2.65 2.645 3.245 ;
      RECT 6.275 2.65 6.605 3.245 ;
      RECT 7.665 2.65 7.995 3.245 ;
      RECT 13.64 2.65 14.23 3.245 ;
      RECT 0.955 2.63 1.205 3.245 ;
      RECT 4.955 2.63 5.205 3.245 ;
  END
END scs8ls_sedfxbp_1

MACRO scs8ls_o32ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.95 3.255 2.12 ;
        RECT 2.925 2.12 3.255 2.735 ;
        RECT 0.565 2.12 0.895 2.735 ;
        RECT 2.925 1.82 3.255 1.95 ;
        RECT 2.925 1.18 3.095 1.82 ;
        RECT 0.545 1.01 3.095 1.18 ;
        RECT 0.545 0.61 0.875 1.01 ;
        RECT 1.545 0.61 1.875 1.01 ;
    END
    ANTENNADIFFAREA 1.1382 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.35 6.115 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.35 4.195 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.35 1.815 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.475 2.905 4.605 3.075 ;
      RECT 4.275 2.29 4.605 2.905 ;
      RECT 3.455 1.95 3.625 2.905 ;
      RECT 2.475 2.29 2.725 2.905 ;
      RECT 3.305 1.01 6.125 1.18 ;
      RECT 3.305 0.84 3.635 1.01 ;
      RECT 4.305 0.35 4.635 1.01 ;
      RECT 5.795 0.35 6.125 1.01 ;
      RECT 2.045 0.67 3.635 0.84 ;
      RECT 2.045 0.425 2.375 0.67 ;
      RECT 3.305 0.35 3.635 0.67 ;
      RECT 0.115 0.255 2.375 0.425 ;
      RECT 0.115 0.425 0.365 1.13 ;
      RECT 1.045 0.425 1.375 0.825 ;
      RECT 0 3.245 6.24 3.415 ;
      RECT 4.835 2.29 5.165 3.245 ;
      RECT 5.87 1.95 6.12 3.245 ;
      RECT 1.465 2.63 1.715 3.245 ;
      RECT 2.555 0.085 3.125 0.5 ;
      RECT 0 -0.085 6.24 0.085 ;
      RECT 3.805 0.085 4.135 0.8 ;
      RECT 4.805 0.085 5.625 0.805 ;
      RECT 0.115 2.905 1.265 3.075 ;
      RECT 1.095 2.46 1.265 2.905 ;
      RECT 1.095 2.29 2.245 2.46 ;
      RECT 1.915 2.46 2.245 2.98 ;
      RECT 0.115 1.95 0.365 2.905 ;
      RECT 3.825 2.12 4.075 2.735 ;
      RECT 3.825 1.95 5.67 2.12 ;
      RECT 5.335 2.12 5.67 2.98 ;
    LAYER mcon ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o32ai_2

MACRO scs8ls_o32ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 11.04 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.765 1.35 10.915 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.35 8.515 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.43 5.635 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.43 4.195 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.43 1.795 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 2.12 1.795 2.735 ;
        RECT 0.645 1.95 5.975 2.12 ;
        RECT 0.645 2.12 0.815 2.735 ;
        RECT 4.735 2.12 5.065 2.735 ;
        RECT 5.635 2.12 5.965 2.735 ;
        RECT 5.805 1.26 5.975 1.95 ;
        RECT 0.545 1.09 5.975 1.26 ;
        RECT 0.545 0.595 0.875 1.09 ;
        RECT 1.555 0.595 1.805 1.09 ;
        RECT 2.475 0.595 2.805 1.09 ;
        RECT 3.475 0.595 3.805 1.09 ;
    END
    ANTENNADIFFAREA 2.2875 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.04 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.04 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.115 2.905 2.245 3.075 ;
      RECT 1.995 2.46 2.245 2.905 ;
      RECT 1.995 2.29 4.055 2.46 ;
      RECT 2.815 2.46 3.145 2.98 ;
      RECT 3.725 2.46 4.055 2.98 ;
      RECT 0.115 1.95 0.445 2.905 ;
      RECT 1.015 2.29 1.265 2.905 ;
      RECT 4.285 2.905 8.465 3.075 ;
      RECT 7.135 2.29 7.465 2.905 ;
      RECT 8.135 2.29 8.465 2.905 ;
      RECT 6.145 1.95 6.465 2.905 ;
      RECT 4.285 2.29 4.535 2.905 ;
      RECT 5.265 2.29 5.435 2.905 ;
      RECT 6.33 1.01 10.67 1.18 ;
      RECT 6.33 0.92 6.67 1.01 ;
      RECT 7.34 0.35 7.67 1.01 ;
      RECT 8.34 0.35 8.67 1.01 ;
      RECT 9.34 0.35 9.67 1.01 ;
      RECT 10.34 0.35 10.67 1.01 ;
      RECT 3.975 0.75 6.67 0.92 ;
      RECT 3.975 0.425 4.305 0.75 ;
      RECT 4.995 0.33 5.325 0.75 ;
      RECT 5.995 0.33 6.67 0.75 ;
      RECT 0.115 0.255 4.305 0.425 ;
      RECT 0.115 0.425 0.365 1.13 ;
      RECT 1.045 0.425 1.375 0.92 ;
      RECT 1.975 0.425 2.305 0.92 ;
      RECT 2.975 0.425 3.305 0.92 ;
      RECT 6.635 2.12 6.965 2.735 ;
      RECT 6.635 1.95 10.475 2.12 ;
      RECT 7.635 2.12 7.965 2.735 ;
      RECT 9.145 2.12 9.475 2.98 ;
      RECT 10.145 2.12 10.475 2.98 ;
      RECT 0 3.245 11.04 3.415 ;
      RECT 8.695 2.29 8.945 3.245 ;
      RECT 9.645 2.29 9.975 3.245 ;
      RECT 10.675 1.95 10.925 3.245 ;
      RECT 2.445 2.63 2.615 3.245 ;
      RECT 3.345 2.63 3.515 3.245 ;
      RECT 4.485 0.085 4.815 0.58 ;
      RECT 0 -0.085 11.04 0.085 ;
      RECT 5.495 0.085 5.825 0.58 ;
      RECT 6.84 0.085 7.17 0.84 ;
      RECT 7.84 0.085 8.17 0.84 ;
      RECT 8.84 0.085 9.17 0.84 ;
      RECT 9.84 0.085 10.17 0.84 ;
    LAYER mcon ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
  END
END scs8ls_o32ai_4

MACRO scs8ls_o41a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.29 0.445 2.98 ;
        RECT 0.115 1.13 0.285 2.29 ;
        RECT 0.115 0.35 0.375 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.3 3.37 2.89 ;
    END
    ANTENNAGATEAREA 0.264 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.47 1.22 2.8 2.89 ;
    END
    ANTENNAGATEAREA 0.264 ;
  END A3

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.61 1.35 4.195 2.15 ;
    END
    ANTENNAGATEAREA 0.264 ;
  END A1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.45 1.58 1.78 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END B1

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.87 1.19 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.264 ;
  END A4

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.875 1.02 4.205 1.03 ;
      RECT 1.675 0.85 4.205 1.02 ;
      RECT 1.675 0.35 2.005 0.85 ;
      RECT 2.675 0.35 3.005 0.85 ;
      RECT 3.875 0.35 4.205 0.85 ;
      RECT 1.75 2.12 2.08 2.845 ;
      RECT 0.455 1.95 2.08 2.12 ;
      RECT 0.615 1.11 1.505 1.28 ;
      RECT 1.175 0.35 1.505 1.11 ;
      RECT 0.455 1.35 0.785 1.95 ;
      RECT 0.615 1.28 0.785 1.35 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 3.76 2.32 4.205 3.245 ;
      RECT 0.615 2.29 1.54 3.245 ;
      RECT 0.545 0.085 0.945 0.94 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 2.175 0.085 2.505 0.68 ;
      RECT 3.175 0.085 3.705 0.68 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o41a_1

MACRO scs8ls_o41a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.95 1.18 4.195 1.41 ;
        RECT 3.95 1.41 4.155 2.98 ;
        RECT 3.95 1.13 4.185 1.18 ;
        RECT 3.855 0.35 4.185 1.13 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.35 3.235 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975 1.35 2.305 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.405 1.35 1.795 1.68 ;
        RECT 1.565 1.68 1.795 2.89 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835 1.92 1.315 2.89 ;
        RECT 0.835 1.35 1.165 1.92 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 0.595 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.115 1.01 2.625 1.18 ;
      RECT 0.115 0.35 0.445 1.01 ;
      RECT 1.115 0.35 1.445 1.01 ;
      RECT 2.295 0.35 2.625 1.01 ;
      RECT 2.125 1.95 3.735 2.12 ;
      RECT 3.405 1.3 3.735 1.95 ;
      RECT 3.405 1.18 3.575 1.3 ;
      RECT 2.795 1.01 3.575 1.18 ;
      RECT 2.795 0.35 3.125 1.01 ;
      RECT 2.125 2.12 2.455 2.98 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 4.355 1.82 4.685 3.245 ;
      RECT 2.695 2.29 3.78 3.245 ;
      RECT 0.115 1.95 0.445 3.245 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 4.355 0.085 4.615 1.01 ;
      RECT 0.615 0.085 0.945 0.84 ;
      RECT 1.615 0.085 2.125 0.815 ;
      RECT 3.355 0.085 3.685 0.82 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o41a_2

MACRO scs8ls_o41a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.425 5.18 1.78 ;
    END
    ANTENNAGATEAREA 0.528 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.875 0.255 4.205 0.67 ;
    END
    ANTENNAGATEAREA 0.528 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805 0.505 8.035 0.67 ;
        RECT 7.305 0.335 8.035 0.505 ;
        RECT 7.305 0.255 7.635 0.335 ;
    END
    ANTENNAGATEAREA 0.528 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.33 1.42 7.075 1.78 ;
    END
    ANTENNAGATEAREA 0.528 ;
  END A1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.94 0.355 2.89 ;
        RECT 0.125 1.77 2.125 1.94 ;
        RECT 0.895 1.94 1.225 2.98 ;
        RECT 1.795 1.94 2.125 2.98 ;
        RECT 0.125 1.1 0.295 1.77 ;
        RECT 0.125 0.93 1.855 1.1 ;
        RECT 0.675 0.35 0.925 0.93 ;
        RECT 1.605 0.35 1.855 0.93 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END X

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.28 1.44 4.195 1.78 ;
    END
    ANTENNAGATEAREA 0.444 ;
  END B1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.455 1.085 7.635 1.25 ;
      RECT 7.385 1.25 7.635 1.275 ;
      RECT 5.665 1.08 7.635 1.085 ;
      RECT 7.385 0.675 7.635 1.08 ;
      RECT 3.455 1.25 5.845 1.255 ;
      RECT 4.725 0.58 4.975 1.085 ;
      RECT 5.665 0.58 5.845 1.08 ;
      RECT 6.455 0.58 6.705 1.08 ;
      RECT 3.455 1.255 3.705 1.27 ;
      RECT 3.455 0.43 3.705 1.085 ;
      RECT 2.595 0.26 3.705 0.43 ;
      RECT 2.595 0.43 2.925 0.93 ;
      RECT 3.79 2.46 4.04 2.98 ;
      RECT 3.79 2.29 5.85 2.46 ;
      RECT 5.68 2.46 5.85 2.98 ;
      RECT 5.68 2.12 5.85 2.29 ;
      RECT 5.68 1.95 7.87 2.12 ;
      RECT 7.54 2.12 7.87 2.98 ;
      RECT 5.68 1.82 5.85 1.95 ;
      RECT 7.54 1.82 7.87 1.95 ;
      RECT 4.24 2.63 5.48 2.98 ;
      RECT 2.78 1.95 5.03 2.12 ;
      RECT 2.78 2.12 3.11 2.79 ;
      RECT 2.78 1.6 3.11 1.95 ;
      RECT 0.585 1.27 3.11 1.6 ;
      RECT 2.94 1.1 3.275 1.27 ;
      RECT 3.105 0.6 3.275 1.1 ;
      RECT 6.05 2.46 6.38 2.98 ;
      RECT 6.05 2.29 7.37 2.46 ;
      RECT 7.04 2.46 7.37 2.98 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 6.58 2.65 6.87 3.245 ;
      RECT 3.31 2.29 3.56 3.245 ;
      RECT 2.325 1.91 2.575 3.245 ;
      RECT 0.525 2.11 0.695 3.245 ;
      RECT 1.425 2.11 1.595 3.245 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 4.375 0.085 4.545 0.915 ;
      RECT 5.155 0.085 5.485 0.915 ;
      RECT 6.025 0.085 6.275 0.91 ;
      RECT 6.885 0.085 7.135 0.91 ;
      RECT 2.035 0.085 2.365 1.1 ;
      RECT 0.175 0.085 0.505 0.76 ;
      RECT 1.105 0.085 1.435 0.76 ;
    LAYER mcon ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
  END
END scs8ls_o41a_4

MACRO scs8ls_o41ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.81 1.35 3.235 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055 1.35 1.385 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A4

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.35 0.775 1.01 ;
        RECT 0.605 1.01 0.775 1.35 ;
        RECT 0.605 1.35 0.885 1.52 ;
        RECT 0.715 1.52 0.885 1.95 ;
        RECT 0.715 1.95 1.165 2.12 ;
        RECT 0.835 2.12 1.165 2.98 ;
    END
    ANTENNADIFFAREA 0.6029 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.435 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.92 2.295 2.89 ;
        RECT 2.125 1.68 2.295 1.92 ;
        RECT 2.125 1.35 2.525 1.68 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.35 1.955 1.68 ;
        RECT 1.565 1.68 1.795 2.89 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A3

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.955 1.01 3.22 1.18 ;
      RECT 0.955 0.35 1.205 1.01 ;
      RECT 1.89 0.35 2.22 1.01 ;
      RECT 2.89 0.35 3.22 1.01 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.995 1.95 3.245 3.245 ;
      RECT 0.115 2.65 0.665 3.245 ;
      RECT 0.115 1.82 0.545 2.65 ;
      RECT 1.375 0.085 1.705 0.84 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.39 0.085 2.72 0.84 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o41ai_1

MACRO scs8ls_o41ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765 1.35 5.155 1.68 ;
        RECT 4.925 1.68 5.155 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.35 3.455 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405 1.35 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A4

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.9 1.55 ;
        RECT 0.125 1.55 0.455 1.63 ;
        RECT 0.125 0.28 0.455 1.18 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 1.55 2.235 1.72 ;
        RECT 0.635 1.72 2.235 1.89 ;
        RECT 1.07 0.645 1.4 1.55 ;
        RECT 0.635 1.89 0.805 2.98 ;
        RECT 2.035 1.89 2.235 2.735 ;
    END
    ANTENNADIFFAREA 0.8792 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.35 1.35 6.115 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 6.24 3.415 ;
      RECT 5.435 2.29 5.605 3.245 ;
      RECT 0.105 1.82 0.435 3.245 ;
      RECT 1.005 2.06 1.335 3.245 ;
      RECT 2.07 0.085 2.4 0.795 ;
      RECT 0 -0.085 6.24 0.085 ;
      RECT 3 0.085 3.33 0.795 ;
      RECT 3.96 0.085 4.29 0.795 ;
      RECT 4.96 0.085 5.29 0.795 ;
      RECT 4.005 2.12 4.335 2.735 ;
      RECT 4.005 1.95 6.135 2.12 ;
      RECT 4.905 2.12 5.235 2.98 ;
      RECT 5.805 2.12 6.135 2.98 ;
      RECT 4.005 1.85 4.335 1.95 ;
      RECT 1.535 2.905 2.765 3.075 ;
      RECT 2.435 2.12 2.765 2.905 ;
      RECT 2.435 1.95 3.8 2.12 ;
      RECT 3.47 2.12 3.8 2.735 ;
      RECT 1.535 2.06 1.865 2.905 ;
      RECT 0.64 0.255 1.9 0.425 ;
      RECT 1.57 0.425 1.9 1.01 ;
      RECT 1.57 1.01 5.79 1.18 ;
      RECT 2.58 0.35 2.83 1.01 ;
      RECT 3.51 0.35 3.79 1.01 ;
      RECT 4.46 0.35 4.79 1.01 ;
      RECT 5.46 0.35 5.79 1.01 ;
      RECT 0.64 0.425 0.89 1.01 ;
      RECT 3.02 2.905 4.705 3.075 ;
      RECT 3.02 2.29 3.27 2.905 ;
      RECT 4.535 2.29 4.705 2.905 ;
    LAYER mcon ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o41ai_2

MACRO scs8ls_o41ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.15 1.89 3.33 2.15 ;
        RECT 2.15 2.15 2.43 2.735 ;
        RECT 3.05 2.15 3.33 2.735 ;
        RECT 0.615 1.72 3.33 1.89 ;
        RECT 0.615 1.89 0.945 2.98 ;
        RECT 1.475 1.01 1.805 1.72 ;
        RECT 0.625 0.84 1.805 1.01 ;
        RECT 0.625 0.595 0.795 0.84 ;
        RECT 1.475 0.595 1.805 0.84 ;
    END
    ANTENNADIFFAREA 1.5862 ;
    ANTENNAPARTIALMETALSIDEAREA 1.389 LAYER li1 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 1.145 1.55 ;
    END
    ANTENNAGATEAREA 0.78 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.142 LAYER li1 ;
  END B1

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.18 3.16 1.55 ;
    END
    ANTENNAGATEAREA 1.116 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.161 LAYER li1 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.395 1.18 6.115 1.55 ;
    END
    ANTENNAGATEAREA 1.116 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.146 LAYER li1 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.18 8.035 1.55 ;
    END
    ANTENNAGATEAREA 1.116 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285 1.18 9.955 1.55 ;
    END
    ANTENNAGATEAREA 1.116 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1 ;
  END A1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.475 0.085 2.99 0.6 ;
      RECT 0 -0.085 10.08 0.085 ;
      RECT 3.67 0.085 3.84 1.13 ;
      RECT 4.52 0.085 4.85 0.67 ;
      RECT 5.45 0.085 5.78 0.67 ;
      RECT 6.38 0.085 6.71 0.67 ;
      RECT 7.24 0.085 7.57 0.67 ;
      RECT 8.205 0.085 8.535 0.67 ;
      RECT 9.205 0.085 9.535 0.67 ;
      RECT 0 3.245 10.08 3.415 ;
      RECT 8.185 2.06 8.515 3.245 ;
      RECT 9.185 2.06 9.515 3.245 ;
      RECT 0.115 1.82 0.445 3.245 ;
      RECT 1.115 2.06 1.445 3.245 ;
      RECT 1.675 2.905 5.705 3.075 ;
      RECT 4.475 2.06 4.805 2.905 ;
      RECT 5.375 2.06 5.705 2.905 ;
      RECT 3.5 1.8 3.805 2.905 ;
      RECT 1.675 2.06 1.98 2.905 ;
      RECT 2.6 2.32 2.88 2.905 ;
      RECT 4.02 0.84 9.965 1.01 ;
      RECT 8.705 0.35 9.035 0.84 ;
      RECT 9.715 0.35 9.965 0.84 ;
      RECT 6.89 0.35 7.06 0.84 ;
      RECT 7.785 0.35 8.035 0.84 ;
      RECT 5.03 0.35 5.28 0.84 ;
      RECT 5.96 0.35 6.21 0.84 ;
      RECT 3.33 1.3 4.19 1.47 ;
      RECT 3.33 1.01 3.5 1.3 ;
      RECT 4.02 1.01 4.19 1.3 ;
      RECT 1.975 0.84 3.5 1.01 ;
      RECT 1.975 0.425 2.305 0.84 ;
      RECT 3.16 0.35 3.5 0.84 ;
      RECT 4.02 0.35 4.35 0.84 ;
      RECT 0.115 0.255 2.305 0.425 ;
      RECT 0.115 0.425 0.445 1.01 ;
      RECT 0.975 0.425 1.305 0.67 ;
      RECT 3.975 1.89 4.305 2.735 ;
      RECT 3.975 1.72 7.565 1.89 ;
      RECT 4.975 1.89 5.205 2.735 ;
      RECT 6.435 1.89 6.665 2.72 ;
      RECT 7.335 1.89 7.565 2.735 ;
      RECT 5.935 2.905 8.015 3.075 ;
      RECT 5.935 2.89 7.165 2.905 ;
      RECT 7.735 1.89 8.015 2.905 ;
      RECT 5.935 2.06 6.265 2.89 ;
      RECT 6.835 2.06 7.165 2.89 ;
      RECT 7.735 1.72 9.965 1.89 ;
      RECT 8.685 1.89 9.015 3 ;
      RECT 9.685 1.89 9.965 3 ;
    LAYER mcon ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o41ai_4

MACRO scs8ls_or2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955 1.82 2.31 2.98 ;
        RECT 2.14 1.13 2.31 1.82 ;
        RECT 1.955 0.35 2.31 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045 1.35 1.375 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.775 1.55 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END B

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.615 1.3 1.97 1.63 ;
      RECT 0.295 1.95 1.785 2.12 ;
      RECT 1.615 1.63 1.785 1.95 ;
      RECT 1.615 1.18 1.785 1.3 ;
      RECT 0.945 1.01 1.785 1.18 ;
      RECT 0.945 0.54 1.24 1.01 ;
      RECT 0.295 2.12 0.625 2.7 ;
      RECT 0.295 1.82 0.625 1.95 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 0.295 0.085 0.65 0.995 ;
      RECT 1.455 0.085 1.785 0.84 ;
      RECT 0 3.245 2.4 3.415 ;
      RECT 1.165 2.29 1.785 3.245 ;
    LAYER mcon ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_or2_1

MACRO scs8ls_or2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.35 1.045 2.15 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.435 1.55 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.555 0.35 1.795 1.82 ;
        RECT 1.555 1.82 1.835 2.15 ;
    END
    ANTENNADIFFAREA 0.5656 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.105 2.32 2.295 2.49 ;
      RECT 2.125 1.63 2.295 2.32 ;
      RECT 1.965 1.3 2.295 1.63 ;
      RECT 1.215 1.18 1.385 2.32 ;
      RECT 0.62 1.01 1.385 1.18 ;
      RECT 0.62 0.45 0.87 1.01 ;
      RECT 0.105 2.49 0.435 2.86 ;
      RECT 0.105 1.82 0.435 2.32 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 1.97 0.085 2.3 1.13 ;
      RECT 0.11 0.085 0.44 1 ;
      RECT 1.045 0.085 1.375 0.825 ;
      RECT 0 3.245 2.4 3.415 ;
      RECT 1.035 2.66 1.365 3.245 ;
      RECT 1.955 2.66 2.285 3.245 ;
    LAYER mcon ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_or2_2

MACRO scs8ls_or2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.21 1.35 2.755 1.95 ;
        RECT 2.52 1.95 3.895 2.12 ;
        RECT 3.59 1.45 3.895 1.95 ;
    END
    ANTENNAGATEAREA 0.411 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.45 3.255 1.78 ;
    END
    ANTENNAGATEAREA 0.411 ;
  END B

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.13 0.355 1.8 ;
        RECT 0.125 1.8 1.795 1.97 ;
        RECT 0.125 0.96 1.7 1.13 ;
        RECT 0.565 1.97 0.895 2.98 ;
        RECT 1.465 1.97 1.795 2.98 ;
        RECT 0.545 0.35 0.795 0.96 ;
        RECT 1.405 0.35 1.7 0.96 ;
    END
    ANTENNADIFFAREA 1.1493 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.45 2.905 3.73 3.075 ;
      RECT 3.4 2.63 3.73 2.905 ;
      RECT 2.45 2.29 2.78 2.905 ;
      RECT 2.98 2.29 4.235 2.46 ;
      RECT 4.065 1.18 4.235 2.29 ;
      RECT 1.87 1.01 4.235 1.18 ;
      RECT 2.98 2.46 3.23 2.735 ;
      RECT 1.87 1.18 2.04 1.3 ;
      RECT 0.595 1.3 2.04 1.63 ;
      RECT 2.42 0.35 2.75 1.01 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 3.93 2.63 4.205 3.245 ;
      RECT 1.995 2.12 2.245 3.245 ;
      RECT 0.115 2.14 0.365 3.245 ;
      RECT 1.095 2.14 1.265 3.245 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 1.92 0.085 2.25 0.84 ;
      RECT 2.92 0.085 4.205 0.84 ;
      RECT 0.115 0.085 0.365 0.79 ;
      RECT 0.975 0.085 1.225 0.79 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_or2_4

MACRO scs8ls_or2b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.035 1.35 2.365 1.78 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END A

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.455 1.55 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END BN

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.755 1.82 3.275 2.98 ;
        RECT 3.105 1.13 3.275 1.82 ;
        RECT 2.875 0.35 3.275 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.115 1.93 0.445 2.98 ;
      RECT 0.115 1.76 0.83 1.93 ;
      RECT 0.66 1.63 0.83 1.76 ;
      RECT 0.66 1.3 1.525 1.63 ;
      RECT 0.66 1.01 0.83 1.3 ;
      RECT 0.115 0.68 0.83 1.01 ;
      RECT 2.535 1.3 2.935 1.63 ;
      RECT 1.695 1.01 2.705 1.18 ;
      RECT 2.535 1.18 2.705 1.3 ;
      RECT 1.695 0.54 2.045 1.01 ;
      RECT 1.3 1.99 1.63 2.86 ;
      RECT 1.3 1.82 1.865 1.99 ;
      RECT 1.695 1.18 1.865 1.82 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 1 0.085 1.525 1.13 ;
      RECT 2.265 0.085 2.68 0.84 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 0.615 2.1 0.945 3.245 ;
      RECT 2.255 1.95 2.585 3.245 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_or2b_1

MACRO scs8ls_or2b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.035 1.35 2.365 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 0.55 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END BN

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.06 0.35 1.39 1.13 ;
        RECT 1.06 1.13 1.23 1.82 ;
        RECT 1.06 1.82 1.645 2.07 ;
    END
    ANTENNADIFFAREA 0.7877 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.875 1.82 3.275 2.86 ;
      RECT 3.105 1.15 3.275 1.82 ;
      RECT 1.625 0.98 3.275 1.15 ;
      RECT 2.405 0.35 2.735 0.98 ;
      RECT 1.625 1.15 1.795 1.3 ;
      RECT 1.465 1.3 1.795 1.63 ;
      RECT 0.115 2.24 2.705 2.41 ;
      RECT 2.535 1.65 2.705 2.24 ;
      RECT 2.535 1.32 2.935 1.65 ;
      RECT 0.115 2.41 0.445 2.7 ;
      RECT 0.115 1.95 0.89 2.24 ;
      RECT 0.72 1.18 0.89 1.95 ;
      RECT 0.12 1.01 0.89 1.18 ;
      RECT 0.12 0.54 0.45 1.01 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 1.56 0.085 2.235 0.81 ;
      RECT 2.915 0.085 3.245 0.81 ;
      RECT 0.63 0.085 0.88 0.84 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 0.65 2.58 0.98 3.245 ;
      RECT 1.765 2.58 2.095 3.245 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_or2b_2

MACRO scs8ls_or2b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.775 1.41 ;
        RECT 0.605 1.41 0.775 1.8 ;
        RECT 0.545 1.13 0.775 1.18 ;
        RECT 0.605 1.8 1.785 1.97 ;
        RECT 0.545 0.96 1.805 1.13 ;
        RECT 0.605 1.97 0.805 2.98 ;
        RECT 1.455 1.97 1.785 2.98 ;
        RECT 0.545 0.35 0.795 0.96 ;
        RECT 1.475 0.35 1.805 0.96 ;
    END
    ANTENNADIFFAREA 1.1049 ;
  END X

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.905 1.12 5.235 1.79 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END BN

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.45 3.235 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.875 1.45 4.125 2.735 ;
      RECT 3.505 1.28 4.125 1.45 ;
      RECT 1.975 1.11 3.755 1.28 ;
      RECT 2.475 0.35 2.805 1.11 ;
      RECT 3.505 0.35 3.755 1.11 ;
      RECT 1.975 1.28 2.145 1.3 ;
      RECT 0.945 1.3 2.145 1.63 ;
      RECT 2.43 2.12 2.76 2.98 ;
      RECT 2.43 1.95 3.675 2.12 ;
      RECT 3.425 2.12 3.675 2.905 ;
      RECT 3.425 1.915 3.675 1.95 ;
      RECT 3.425 2.905 4.655 3.075 ;
      RECT 4.325 1.945 4.655 2.905 ;
      RECT 4.435 0.35 5.655 0.95 ;
      RECT 5.405 0.95 5.655 2.98 ;
      RECT 4.295 1.445 4.625 1.775 ;
      RECT 4.435 0.95 4.625 1.445 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 2.96 2.29 3.21 3.245 ;
      RECT 4.875 1.96 5.205 3.245 ;
      RECT 1.985 1.94 2.235 3.245 ;
      RECT 0.105 1.82 0.435 3.245 ;
      RECT 1.005 2.14 1.255 3.245 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 1.975 0.085 2.305 0.94 ;
      RECT 3.005 0.085 3.335 0.94 ;
      RECT 3.935 0.085 4.265 1.03 ;
      RECT 0.115 0.085 0.365 1.01 ;
      RECT 0.975 0.085 1.305 0.765 ;
    LAYER mcon ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_or2b_4

MACRO scs8ls_or3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.43 0.35 2.795 1.13 ;
        RECT 2.625 1.13 2.795 1.82 ;
        RECT 2.515 1.82 2.795 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 0.57 1.78 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835 1.35 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.35 1.815 1.78 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.09 1.3 2.455 1.63 ;
      RECT 0.115 1.95 2.26 2.12 ;
      RECT 2.09 1.63 2.26 1.95 ;
      RECT 2.09 1.18 2.26 1.3 ;
      RECT 0.115 1.01 2.26 1.18 ;
      RECT 1.045 0.455 1.76 1.01 ;
      RECT 0.115 2.12 0.445 2.86 ;
      RECT 0.115 0.35 0.365 1.01 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 1.555 2.29 2.315 3.245 ;
      RECT 0 -0.085 2.88 0.085 ;
      RECT 0.545 0.085 0.875 0.81 ;
      RECT 1.93 0.085 2.26 0.81 ;
    LAYER mcon ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
  END
END scs8ls_or3_1

MACRO scs8ls_or3_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.13 1.335 2.89 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.18 1.905 1.55 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.12 0.835 1.79 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END C

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.13 3.235 1.8 ;
        RECT 2.335 1.8 3.235 1.97 ;
        RECT 2.415 0.96 3.235 1.13 ;
        RECT 2.335 1.97 2.665 2.98 ;
        RECT 2.415 0.35 2.745 0.96 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.075 1.3 2.815 1.63 ;
      RECT 0.095 0.79 2.245 0.95 ;
      RECT 1.2 0.95 2.245 0.96 ;
      RECT 2.075 0.96 2.245 1.3 ;
      RECT 0.095 0.78 1.53 0.79 ;
      RECT 1.2 0.35 1.53 0.78 ;
      RECT 0.285 2.13 0.615 2.98 ;
      RECT 0.095 1.96 0.615 2.13 ;
      RECT 0.095 0.35 0.445 0.78 ;
      RECT 0.095 0.95 0.265 1.96 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.835 2.14 3.165 3.245 ;
      RECT 1.725 1.94 2.055 3.245 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.915 0.085 3.245 0.79 ;
      RECT 0.615 0.085 1.03 0.6 ;
      RECT 1.7 0.085 2.245 0.6 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_or3_2

MACRO scs8ls_or3_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.13 5.155 1.8 ;
        RECT 3.565 1.8 5.155 1.97 ;
        RECT 3.565 0.96 5.155 1.13 ;
        RECT 3.565 1.97 3.735 2.98 ;
        RECT 4.385 1.97 4.715 2.98 ;
        RECT 3.565 0.35 3.735 0.96 ;
        RECT 4.405 0.35 4.655 0.96 ;
    END
    ANTENNADIFFAREA 1.0901 ;
  END X

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.05 0.27 1.38 0.94 ;
    END
    ANTENNAGATEAREA 0.411 ;
  END C

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.28 0.435 1.63 ;
        RECT 0.105 1.11 3.055 1.28 ;
        RECT 2.755 1.28 3.055 1.55 ;
        RECT 0.105 0.28 0.435 1.11 ;
    END
    ANTENNAGATEAREA 0.411 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.45 2.545 1.78 ;
    END
    ANTENNAGATEAREA 0.411 ;
  END B

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.28 0.085 ;
      RECT 4.835 0.085 5.165 0.79 ;
      RECT 2.05 0.085 2.38 0.6 ;
      RECT 3.05 0.085 3.38 0.6 ;
      RECT 3.915 0.085 4.165 0.79 ;
      RECT 1.015 2.71 2.33 2.96 ;
      RECT 3.225 1.3 4.685 1.63 ;
      RECT 1.495 1.95 3.395 2.12 ;
      RECT 3.225 1.63 3.395 1.95 ;
      RECT 3.225 0.94 3.395 1.3 ;
      RECT 1.55 0.77 3.395 0.94 ;
      RECT 2.55 0.35 2.88 0.77 ;
      RECT 1.495 2.12 1.825 2.2 ;
      RECT 1.55 0.35 1.88 0.77 ;
      RECT 0.565 2.54 0.815 2.96 ;
      RECT 0.565 2.37 2.83 2.54 ;
      RECT 2.5 2.54 2.83 2.96 ;
      RECT 2.5 2.29 2.83 2.37 ;
      RECT 0.565 1.95 0.815 2.37 ;
      RECT 0 3.245 5.28 3.415 ;
      RECT 4.915 2.14 5.165 3.245 ;
      RECT 3.035 2.29 3.365 3.245 ;
      RECT 0.115 1.92 0.365 3.245 ;
      RECT 3.935 2.14 4.185 3.245 ;
    LAYER mcon ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_or3_4

MACRO scs8ls_or3b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395 0.35 3.755 1.13 ;
        RECT 3.585 1.13 3.755 1.82 ;
        RECT 3.25 1.82 3.755 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.11 0.605 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END CN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.915 1.19 2.275 2.89 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.515 1.3 2.845 1.78 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.615 2.1 0.945 2.98 ;
      RECT 0.775 1.88 0.945 2.1 ;
      RECT 0.775 1.21 1.205 1.88 ;
      RECT 0.775 0.94 0.945 1.21 ;
      RECT 0.615 0.35 0.945 0.94 ;
      RECT 3.055 1.3 3.415 1.63 ;
      RECT 3.055 1.02 3.225 1.3 ;
      RECT 1.175 0.85 3.225 1.02 ;
      RECT 2.175 0.35 2.505 0.85 ;
      RECT 1.375 1.02 1.705 2.975 ;
      RECT 1.175 0.35 1.505 0.85 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 2.75 1.95 3.08 3.245 ;
      RECT 0.115 2.1 0.445 3.245 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 0.115 0.085 0.445 0.94 ;
      RECT 1.675 0.085 2.005 0.68 ;
      RECT 2.675 0.085 3.225 0.68 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_or3b_1

MACRO scs8ls_or3b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.3 0.435 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END CN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.515 1.35 2.845 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975 1.35 2.305 2.15 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.82 1.795 2.15 ;
        RECT 1.065 1.13 1.235 1.82 ;
        RECT 1.065 0.96 1.455 1.13 ;
        RECT 1.125 0.35 1.455 0.96 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.115 2.32 2.645 2.49 ;
      RECT 2.475 2.12 2.645 2.32 ;
      RECT 2.475 1.95 3.415 2.12 ;
      RECT 3.085 1.35 3.415 1.95 ;
      RECT 0.115 2.49 0.445 2.7 ;
      RECT 0.115 1.95 0.775 2.32 ;
      RECT 0.605 1.13 0.775 1.95 ;
      RECT 0.185 0.96 0.775 1.13 ;
      RECT 0.185 0.54 0.605 0.96 ;
      RECT 3.235 2.29 3.755 2.86 ;
      RECT 3.585 1.18 3.755 2.29 ;
      RECT 1.625 1.01 3.755 1.18 ;
      RECT 2.35 0.45 2.68 1.01 ;
      RECT 3.35 0.45 3.755 1.01 ;
      RECT 1.625 1.18 1.795 1.3 ;
      RECT 1.405 1.3 1.795 1.63 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 0.65 2.66 0.98 3.245 ;
      RECT 1.635 2.66 2.07 3.245 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 1.625 0.085 2.135 0.78 ;
      RECT 2.85 0.085 3.18 0.84 ;
      RECT 0.775 0.085 0.945 0.79 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_or3b_2

MACRO scs8ls_or3b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405 1.13 5.635 1.8 ;
        RECT 4.055 1.8 5.635 1.97 ;
        RECT 4.055 0.96 5.635 1.13 ;
        RECT 4.055 1.97 4.225 2.98 ;
        RECT 4.875 1.97 5.205 2.98 ;
        RECT 4.055 0.35 4.225 0.96 ;
        RECT 4.885 0.35 5.135 0.96 ;
    END
    ANTENNADIFFAREA 1.1049 ;
  END X

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.255 0.775 0.64 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END CN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.34 1.55 3.075 1.8 ;
        RECT 1.34 1.49 1.67 1.55 ;
    END
    ANTENNAGATEAREA 0.411 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.8 1.15 3.545 1.32 ;
        RECT 3.005 1.32 3.545 1.38 ;
        RECT 0.8 1.32 1.13 1.76 ;
        RECT 3.285 1.38 3.545 1.55 ;
    END
    ANTENNAGATEAREA 0.411 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 5.405 2.14 5.655 3.245 ;
      RECT 3.505 2.31 3.835 3.245 ;
      RECT 0.56 1.94 0.89 3.245 ;
      RECT 4.425 2.14 4.675 3.245 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 5.315 0.085 5.645 0.79 ;
      RECT 0.945 0.085 1.41 0.64 ;
      RECT 2.58 0.085 2.91 0.64 ;
      RECT 3.51 0.085 3.85 0.6 ;
      RECT 4.405 0.085 4.655 0.79 ;
      RECT 1.58 2.7 2.835 2.98 ;
      RECT 0.11 0.81 1.91 0.98 ;
      RECT 1.58 0.31 1.91 0.81 ;
      RECT 0.11 1.34 0.36 2.98 ;
      RECT 0.11 0.98 0.465 1.34 ;
      RECT 3.715 1.3 5.175 1.63 ;
      RECT 2.03 1.97 3.885 2.14 ;
      RECT 3.715 1.63 3.885 1.97 ;
      RECT 3.715 0.98 3.885 1.3 ;
      RECT 2.08 0.81 3.885 0.98 ;
      RECT 3.09 0.35 3.34 0.81 ;
      RECT 2.03 2.14 2.385 2.19 ;
      RECT 2.08 0.35 2.41 0.81 ;
      RECT 1.07 2.53 1.4 2.98 ;
      RECT 1.07 2.36 3.335 2.53 ;
      RECT 3.005 2.53 3.335 2.98 ;
      RECT 3.005 2.31 3.335 2.36 ;
      RECT 1.07 1.97 1.4 2.36 ;
    LAYER mcon ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_or3b_4

MACRO scs8ls_or4_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.49 1.42 1.82 1.78 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END B

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.9 1.82 3.275 2.98 ;
        RECT 3.105 1.13 3.275 1.82 ;
        RECT 2.96 0.35 3.275 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 2.39 1.78 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.92 1.42 1.295 1.78 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.42 0.65 1.78 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.56 1.3 2.935 1.63 ;
      RECT 0.2 1.95 2.73 2.12 ;
      RECT 2.56 1.63 2.73 1.95 ;
      RECT 2.56 1.18 2.73 1.3 ;
      RECT 0.615 1.01 2.73 1.18 ;
      RECT 1.86 0.54 2.19 1.01 ;
      RECT 0.615 0.54 0.945 1.01 ;
      RECT 0.2 2.12 0.53 2.98 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 0.115 0.085 0.445 1.13 ;
      RECT 1.125 0.085 1.6 0.84 ;
      RECT 2.45 0.085 2.78 0.84 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.15 2.29 2.565 3.245 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_or4_1

MACRO scs8ls_or4_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.165 1.335 2.89 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.35 1.875 2.89 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 2.455 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.18 0.835 1.77 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END D

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.13 3.715 1.8 ;
        RECT 2.86 1.8 3.715 1.97 ;
        RECT 2.965 0.96 3.715 1.13 ;
        RECT 2.86 1.97 3.19 2.98 ;
        RECT 2.965 0.35 3.215 0.96 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.625 1.3 3.04 1.63 ;
      RECT 0.085 0.825 2.19 0.995 ;
      RECT 1.86 0.995 2.19 1.01 ;
      RECT 1.86 0.35 2.19 0.825 ;
      RECT 1.86 1.01 2.795 1.18 ;
      RECT 2.625 1.18 2.795 1.3 ;
      RECT 0.69 0.35 1.02 0.825 ;
      RECT 0.405 2.11 0.735 2.98 ;
      RECT 0.085 1.94 0.735 2.11 ;
      RECT 0.085 0.995 0.255 1.94 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 3.36 2.14 3.69 3.245 ;
      RECT 2.36 1.95 2.69 3.245 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 3.395 0.085 3.725 0.775 ;
      RECT 0.115 0.085 0.51 0.655 ;
      RECT 1.2 0.085 1.68 0.655 ;
      RECT 2.36 0.085 2.795 0.825 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_or4_2

MACRO scs8ls_or4_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.47 3.735 1.8 ;
    END
    ANTENNAGATEAREA 0.411 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.13 4.395 1.3 ;
        RECT 2.525 1.3 3.235 1.41 ;
        RECT 4.065 1.3 4.395 1.55 ;
        RECT 2.615 1.41 3.235 1.55 ;
    END
    ANTENNAGATEAREA 0.411 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.605 1.365 6.285 1.77 ;
        RECT 4.925 1.77 6.285 1.78 ;
    END
    ANTENNAGATEAREA 0.411 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.285 0.255 6.615 0.855 ;
    END
    ANTENNAGATEAREA 0.411 ;
  END D

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.82 2.275 2.15 ;
        RECT 0.615 2.15 0.845 2.98 ;
        RECT 1.515 2.15 1.745 2.98 ;
        RECT 0.125 1.3 0.945 1.82 ;
        RECT 0.615 1.15 0.945 1.3 ;
        RECT 0.615 0.98 1.945 1.15 ;
        RECT 0.615 0.35 0.945 0.98 ;
        RECT 1.615 0.35 1.945 0.98 ;
    END
    ANTENNADIFFAREA 1.3269 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.72 0.085 ;
      RECT 2.38 0.085 2.74 0.62 ;
      RECT 3.43 0.085 4.59 0.62 ;
      RECT 5.27 0.085 6.115 0.68 ;
      RECT 0.115 0.085 0.445 1.13 ;
      RECT 1.115 0.085 1.445 0.81 ;
      RECT 0 3.245 6.72 3.415 ;
      RECT 3.375 2.73 3.705 3.245 ;
      RECT 1.915 2.32 2.245 3.245 ;
      RECT 0.115 2.32 0.445 3.245 ;
      RECT 1.015 2.32 1.345 3.245 ;
      RECT 5.295 1.95 6.635 2.12 ;
      RECT 6.465 1.195 6.635 1.95 ;
      RECT 4.77 1.025 6.635 1.195 ;
      RECT 5.295 2.12 5.625 2.19 ;
      RECT 4.77 0.96 5.1 1.025 ;
      RECT 2.155 0.79 5.1 0.96 ;
      RECT 4.77 0.35 5.1 0.79 ;
      RECT 2.155 0.96 2.325 1.32 ;
      RECT 1.315 1.32 2.325 1.65 ;
      RECT 2.92 0.35 3.25 0.79 ;
      RECT 4.345 2.53 4.675 2.98 ;
      RECT 4.345 2.36 6.575 2.53 ;
      RECT 6.245 2.53 6.575 2.98 ;
      RECT 6.245 2.29 6.575 2.36 ;
      RECT 4.345 2.14 4.675 2.36 ;
      RECT 2.475 1.97 4.675 2.14 ;
      RECT 2.475 2.14 2.805 2.19 ;
      RECT 2.475 1.94 2.805 1.97 ;
      RECT 4.345 1.94 4.675 1.97 ;
      RECT 2.475 2.19 2.755 2.98 ;
      RECT 4.845 2.7 6.075 2.98 ;
      RECT 2.925 2.56 3.205 2.98 ;
      RECT 2.925 2.36 4.175 2.56 ;
      RECT 3.895 2.56 4.175 2.98 ;
      RECT 3.825 2.31 4.175 2.36 ;
    LAYER mcon ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_or4_4

MACRO scs8ls_or4b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.835 1.82 4.235 2.98 ;
        RECT 4.065 1.13 4.235 1.82 ;
        RECT 3.835 0.35 4.235 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885 1.045 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.455 1.18 2.785 1.78 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.995 1.35 3.325 1.78 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END A

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.45 0.57 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END DN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.495 1.3 3.895 1.63 ;
      RECT 1.315 1.95 3.665 2.12 ;
      RECT 3.495 1.63 3.665 1.95 ;
      RECT 3.495 1.18 3.665 1.3 ;
      RECT 2.955 1.01 3.665 1.18 ;
      RECT 2.955 0.94 3.125 1.01 ;
      RECT 2.76 0.35 3.125 0.94 ;
      RECT 1.115 0.545 2.09 0.875 ;
      RECT 1.315 2.12 1.645 2.86 ;
      RECT 1.315 0.875 1.645 1.95 ;
      RECT 0.12 2.12 0.45 2.98 ;
      RECT 0.12 1.95 0.98 2.12 ;
      RECT 0.81 1.91 0.98 1.95 ;
      RECT 0.81 1.58 1.14 1.91 ;
      RECT 0.81 1.28 0.98 1.58 ;
      RECT 0.115 1.11 0.98 1.28 ;
      RECT 0.115 0.35 0.445 1.11 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 0.62 2.29 0.95 3.245 ;
      RECT 3.335 2.29 3.665 3.245 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 0.615 0.085 0.945 0.94 ;
      RECT 2.26 0.085 2.59 0.875 ;
      RECT 3.295 0.085 3.625 0.84 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_or4b_1

MACRO scs8ls_or4b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.06 1.82 1.43 2.15 ;
        RECT 1.06 1.13 1.23 1.82 ;
        RECT 1.06 0.35 1.405 1.13 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 0.55 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END DN

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.47 3.355 2.52 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.485 1.47 2.815 2.15 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945 1.35 2.275 2.15 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.865 1.94 4.235 2.98 ;
      RECT 4.065 1.27 4.235 1.94 ;
      RECT 3.375 1.13 4.235 1.27 ;
      RECT 1.575 1.1 4.235 1.13 ;
      RECT 1.575 0.96 3.705 1.1 ;
      RECT 3.375 0.45 3.705 0.96 ;
      RECT 2.175 0.45 2.505 0.96 ;
      RECT 1.575 1.13 1.745 1.3 ;
      RECT 1.4 1.3 1.745 1.63 ;
      RECT 2.295 2.69 3.695 2.86 ;
      RECT 3.525 1.77 3.695 2.69 ;
      RECT 3.525 1.44 3.895 1.77 ;
      RECT 0.115 2.32 2.465 2.49 ;
      RECT 2.295 2.49 2.465 2.69 ;
      RECT 0.115 2.49 0.445 2.7 ;
      RECT 0.115 1.95 0.89 2.32 ;
      RECT 0.72 1.18 0.89 1.95 ;
      RECT 0.13 1.01 0.89 1.18 ;
      RECT 0.13 0.54 0.46 1.01 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 1.55 2.73 2.125 3.245 ;
      RECT 0.65 2.66 0.98 3.245 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 1.575 0.085 1.995 0.78 ;
      RECT 2.685 0.085 3.205 0.78 ;
      RECT 3.875 0.085 4.205 0.93 ;
      RECT 0.64 0.085 0.89 0.84 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_or4b_2

MACRO scs8ls_or4b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.18 4.815 1.55 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END DN

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.41 1.82 7.075 2.15 ;
        RECT 5.41 2.15 5.69 2.98 ;
        RECT 6.365 1.47 6.655 1.82 ;
        RECT 6.325 1.3 6.655 1.47 ;
        RECT 6.325 1.15 6.575 1.3 ;
        RECT 5.325 0.98 6.575 1.15 ;
        RECT 5.325 0.35 5.655 0.98 ;
        RECT 6.325 0.35 6.575 0.98 ;
        RECT 6.36 2.15 6.59 2.98 ;
    END
    ANTENNADIFFAREA 1.1789 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.45 1.335 1.78 ;
    END
    ANTENNAGATEAREA 0.411 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.28 0.835 1.55 ;
        RECT 0.125 1.11 2.035 1.28 ;
        RECT 1.705 1.28 2.035 1.55 ;
    END
    ANTENNAGATEAREA 0.411 ;
  END B

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
    END
  END vpwr

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2.495 1.225 4.225 1.365 ;
        RECT 2.495 1.365 2.785 1.41 ;
        RECT 2.495 1.18 2.785 1.225 ;
        RECT 3.935 1.365 4.225 1.41 ;
        RECT 3.935 1.18 4.225 1.225 ;
    END
    ANTENNAGATEAREA 0.411 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.197 LAYER met1 ;
  END C

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.245 1.18 2.725 1.78 ;
      RECT 3.865 1.18 4.195 1.51 ;
      RECT 0.645 2.46 0.815 2.98 ;
      RECT 0.645 2.29 1.845 2.46 ;
      RECT 1.515 2.46 1.845 2.98 ;
      RECT 2.015 2.53 2.345 2.98 ;
      RECT 2.015 2.36 4.195 2.53 ;
      RECT 3.945 2.53 4.195 2.98 ;
      RECT 2.015 2.12 2.345 2.36 ;
      RECT 3.945 2.06 4.195 2.36 ;
      RECT 0.115 1.95 2.345 2.12 ;
      RECT 0.115 2.12 0.445 2.98 ;
      RECT 0.115 1.94 0.445 1.95 ;
      RECT 2.515 2.7 3.745 2.98 ;
      RECT 3.44 0.34 4.565 0.67 ;
      RECT 4.425 1.89 4.755 2.86 ;
      RECT 3.465 1.8 4.755 1.89 ;
      RECT 3.235 1.72 4.755 1.8 ;
      RECT 3.235 1.47 3.635 1.72 ;
      RECT 4.985 1.32 6.155 1.65 ;
      RECT 2.895 0.94 5.155 1.01 ;
      RECT 4.985 1.01 5.155 1.32 ;
      RECT 0.115 0.84 5.155 0.94 ;
      RECT 2.895 2.02 3.295 2.19 ;
      RECT 2.895 1.13 3.065 2.02 ;
      RECT 2.895 1.01 3.27 1.13 ;
      RECT 0.115 0.77 3.27 0.84 ;
      RECT 1.115 0.35 2.2 0.77 ;
      RECT 2.895 0.35 3.27 0.77 ;
      RECT 0.115 0.35 0.445 0.77 ;
      RECT 0 -0.085 7.2 0.085 ;
      RECT 6.755 0.085 7.085 1.13 ;
      RECT 0.615 0.085 0.945 0.6 ;
      RECT 2.37 0.085 2.725 0.6 ;
      RECT 4.825 0.085 5.155 0.67 ;
      RECT 5.825 0.085 6.155 0.81 ;
      RECT 0 3.245 7.2 3.415 ;
      RECT 6.76 2.32 7.09 3.245 ;
      RECT 1.015 2.63 1.345 3.245 ;
      RECT 4.96 1.82 5.21 3.245 ;
      RECT 5.86 2.32 6.19 3.245 ;
    LAYER mcon ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.555 1.21 2.725 1.38 ;
      RECT 3.995 1.21 4.165 1.38 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
  END
END scs8ls_or4b_4

MACRO scs8ls_o22a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.45 3.505 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B2

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.845 1.45 1.515 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.845 1.45 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.935 1.18 6.595 1.41 ;
        RECT 5.935 1.41 6.105 1.85 ;
        RECT 4.98 1.01 6.105 1.18 ;
        RECT 4.6 1.85 6.105 2.02 ;
        RECT 4.98 0.35 5.23 1.01 ;
        RECT 5.92 0.35 6.105 1.01 ;
        RECT 4.6 2.02 4.93 2.98 ;
        RECT 5.775 2.02 6.105 2.98 ;
    END
    ANTENNADIFFAREA 1.1256 ;
  END X

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 0.255 2.61 0.57 ;
        RECT 2.045 0.57 2.275 0.67 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.565 2.905 3.895 3.075 ;
      RECT 2.565 2.29 2.895 2.905 ;
      RECT 3.565 2.29 3.895 2.905 ;
      RECT 0 3.245 6.72 3.415 ;
      RECT 6.275 1.82 6.605 3.245 ;
      RECT 2.065 2.29 2.395 3.245 ;
      RECT 0.115 1.94 0.365 3.245 ;
      RECT 4.1 1.85 4.43 3.245 ;
      RECT 5.2 2.19 5.53 3.245 ;
      RECT 0 -0.085 6.72 0.085 ;
      RECT 6.275 0.085 6.605 1.01 ;
      RECT 4.47 0.085 4.8 0.58 ;
      RECT 5.41 0.085 5.74 0.79 ;
      RECT 0.615 0.085 0.945 0.94 ;
      RECT 1.545 0.085 1.875 0.94 ;
      RECT 3.675 1.51 5.765 1.68 ;
      RECT 4.415 1.35 5.765 1.51 ;
      RECT 1.065 1.95 3.845 2.12 ;
      RECT 3.065 2.12 3.395 2.735 ;
      RECT 3.675 1.68 3.845 1.95 ;
      RECT 4.415 0.92 4.585 1.35 ;
      RECT 2.545 0.75 4.585 0.92 ;
      RECT 2.545 0.74 3.81 0.75 ;
      RECT 3.48 0.66 3.81 0.74 ;
      RECT 1.065 2.12 1.395 2.735 ;
      RECT 0.115 1.11 4.24 1.28 ;
      RECT 3.91 1.28 4.24 1.34 ;
      RECT 2.045 1.09 4.24 1.11 ;
      RECT 2.045 0.84 2.375 1.09 ;
      RECT 0.115 1.28 0.445 1.34 ;
      RECT 0.115 0.66 0.445 1.11 ;
      RECT 1.125 0.66 1.375 1.11 ;
      RECT 0.565 2.905 1.895 3.075 ;
      RECT 1.565 2.29 1.895 2.905 ;
      RECT 0.565 1.95 0.895 2.905 ;
    LAYER mcon ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o22a_4

MACRO scs8ls_o22ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.3 2.775 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535 1.35 1.865 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625 1.95 1.55 2.98 ;
        RECT 0.625 1.13 0.795 1.95 ;
        RECT 0.615 0.655 1.065 1.13 ;
    END
    ANTENNADIFFAREA 0.8959 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.18 0.445 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.35 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.115 0.315 1.67 0.485 ;
      RECT 1.34 0.485 1.67 0.96 ;
      RECT 1.34 0.96 2.67 1.13 ;
      RECT 2.34 0.35 2.67 0.96 ;
      RECT 0.115 0.485 0.445 1.01 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 2.255 1.95 2.585 3.245 ;
      RECT 0.125 1.82 0.455 3.245 ;
      RECT 1.84 0.085 2.17 0.79 ;
      RECT 0 -0.085 2.88 0.085 ;
    LAYER mcon ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o22ai_1

MACRO scs8ls_o22ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.18 2.275 1.8 ;
        RECT 2.045 1.8 3.31 1.95 ;
        RECT 0.615 1.01 2.275 1.18 ;
        RECT 1.57 1.95 3.31 1.97 ;
        RECT 0.615 0.595 0.945 1.01 ;
        RECT 1.615 0.595 1.945 1.01 ;
        RECT 1.57 1.97 2.275 2.12 ;
        RECT 3.06 1.97 3.31 2.735 ;
        RECT 1.57 2.12 1.8 2.735 ;
    END
    ANTENNADIFFAREA 1.2122 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.91 1.35 4.675 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.63 3.715 1.78 ;
        RECT 2.665 1.39 3.715 1.63 ;
        RECT 2.665 1.3 3.335 1.39 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.35 1.815 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.53 2.905 3.68 3.075 ;
      RECT 3.51 2.12 3.68 2.905 ;
      RECT 3.51 1.95 4.66 2.12 ;
      RECT 4.33 2.12 4.66 2.98 ;
      RECT 2.53 2.14 2.86 2.905 ;
      RECT 1.07 2.905 2.3 3.075 ;
      RECT 1.97 2.29 2.3 2.905 ;
      RECT 1.07 2.12 1.4 2.905 ;
      RECT 0.12 1.95 1.4 2.12 ;
      RECT 0.12 2.12 0.37 2.98 ;
      RECT 3.505 1.13 4.685 1.18 ;
      RECT 2.455 1.01 4.685 1.13 ;
      RECT 2.455 0.96 3.755 1.01 ;
      RECT 4.435 0.35 4.685 1.01 ;
      RECT 2.455 0.84 2.785 0.96 ;
      RECT 3.505 0.35 3.755 0.96 ;
      RECT 2.115 0.425 2.785 0.84 ;
      RECT 0.115 0.255 2.785 0.425 ;
      RECT 0.115 0.425 0.445 1.13 ;
      RECT 1.115 0.425 1.445 0.84 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 3.88 2.29 4.13 3.245 ;
      RECT 0.57 2.29 0.9 3.245 ;
      RECT 2.955 0.085 3.285 0.79 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 3.925 0.085 4.255 0.84 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o22ai_2

MACRO scs8ls_o22ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.89 3.235 2.15 ;
        RECT 1.38 1.72 3.81 1.89 ;
        RECT 3.64 1.68 3.81 1.72 ;
        RECT 1.38 1.65 1.55 1.72 ;
        RECT 3.64 1.35 3.97 1.68 ;
        RECT 0.54 1.32 1.55 1.65 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885 1.18 3.235 1.55 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.405 0.92 5.155 1.13 ;
        RECT 4.405 0.75 8.07 0.92 ;
        RECT 7.9 0.92 8.07 1.95 ;
        RECT 6.205 0.595 6.535 0.75 ;
        RECT 7.205 0.595 7.535 0.75 ;
        RECT 3.98 1.95 8.07 2.02 ;
        RECT 3.98 2.02 4.15 2.32 ;
        RECT 5.77 2.02 8.07 2.12 ;
        RECT 3.98 1.85 6.1 1.95 ;
        RECT 2.02 2.32 4.15 2.49 ;
        RECT 5.77 2.12 6.1 2.735 ;
        RECT 6.67 2.12 7 2.735 ;
        RECT 2.02 2.06 2.35 2.32 ;
    END
    ANTENNADIFFAREA 2.388 ;
  END Y

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.805 1.43 7.155 1.68 ;
        RECT 6.365 1.68 7.155 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405 1.26 5.635 1.3 ;
        RECT 4.29 1.3 5.635 1.63 ;
        RECT 5.405 1.09 7.73 1.26 ;
        RECT 7.4 1.26 7.73 1.55 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.905 0.255 8.045 0.425 ;
      RECT 7.715 0.425 8.045 0.58 ;
      RECT 3.905 0.425 6.035 0.58 ;
      RECT 6.705 0.425 7.035 0.58 ;
      RECT 0.115 1.01 1.375 1.15 ;
      RECT 0.115 0.98 4.235 1.01 ;
      RECT 3.905 1.01 4.235 1.13 ;
      RECT 1.125 0.84 4.235 0.98 ;
      RECT 0.115 0.35 0.445 0.98 ;
      RECT 3.905 0.58 4.235 0.84 ;
      RECT 1.125 0.35 1.375 0.84 ;
      RECT 2.055 0.35 2.305 0.84 ;
      RECT 2.985 0.35 3.235 0.84 ;
      RECT 5.32 2.905 7.5 3.075 ;
      RECT 7.17 2.29 7.5 2.905 ;
      RECT 4.37 2.36 4.7 2.98 ;
      RECT 4.37 2.19 5.57 2.36 ;
      RECT 5.32 2.36 5.57 2.905 ;
      RECT 6.3 2.29 6.47 2.905 ;
      RECT 1.52 2.66 3.7 2.98 ;
      RECT 0.57 2.23 0.85 2.98 ;
      RECT 0.57 1.82 0.9 2.06 ;
      RECT 1.52 2.23 1.85 2.66 ;
      RECT 0.57 2.06 1.85 2.23 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 7.67 2.29 8 3.245 ;
      RECT 1.02 2.4 1.35 3.245 ;
      RECT 0.12 1.82 0.37 3.245 ;
      RECT 3.87 2.66 4.2 3.245 ;
      RECT 4.9 2.53 5.15 3.245 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 0.615 0.085 0.945 0.81 ;
      RECT 1.545 0.085 1.875 0.67 ;
      RECT 2.475 0.085 2.805 0.67 ;
      RECT 3.405 0.085 3.735 0.67 ;
    LAYER mcon ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
  END
END scs8ls_o22ai_4

MACRO scs8ls_o2bb2a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.42 1.315 1.71 ;
        RECT 1.085 1.71 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END A1N

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885 1.18 4.215 1.51 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.82 0.445 2.98 ;
        RECT 0.085 1.13 0.255 1.82 ;
        RECT 0.085 0.35 0.455 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.43 1.835 1.78 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END A2N

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.18 3.715 1.51 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.15 1.95 2.38 2.28 ;
      RECT 2.05 1.26 2.38 1.95 ;
      RECT 1.63 1.09 2.38 1.26 ;
      RECT 1.63 0.595 1.88 1.09 ;
      RECT 2.995 0.84 4.205 1.01 ;
      RECT 2.995 0.34 3.245 0.84 ;
      RECT 3.955 0.34 4.205 0.84 ;
      RECT 2.99 2.07 3.32 2.78 ;
      RECT 2.645 1.9 3.32 2.07 ;
      RECT 2.645 0.92 2.815 1.9 ;
      RECT 2.485 0.425 2.815 0.92 ;
      RECT 1.29 0.255 2.815 0.425 ;
      RECT 1.29 0.425 1.46 1.08 ;
      RECT 0.625 1.08 1.46 1.25 ;
      RECT 0.625 1.25 0.795 1.3 ;
      RECT 0.425 1.3 0.795 1.63 ;
      RECT 0.625 0.085 1.12 0.91 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 3.415 0.085 3.745 0.67 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 1.655 2.45 2.82 3.245 ;
      RECT 0.615 1.95 0.945 3.245 ;
      RECT 3.87 1.9 4.2 3.245 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_o2bb2a_1

MACRO scs8ls_o2bb2a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.81 1.45 1.285 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.45 0.57 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.425 1.82 3.77 2.98 ;
        RECT 3.6 1.13 3.77 1.82 ;
        RECT 3.43 0.35 3.77 1.13 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.995 1.475 2.325 1.805 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END A2N

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.475 2.865 1.805 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END A1N

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.085 1.305 3.43 1.635 ;
      RECT 1.05 2.395 3.255 2.565 ;
      RECT 3.085 1.635 3.255 2.395 ;
      RECT 2.545 1.135 3.255 1.305 ;
      RECT 2.545 0.425 2.715 1.135 ;
      RECT 1.475 0.255 2.715 0.425 ;
      RECT 1.05 2.565 1.38 2.98 ;
      RECT 1.05 1.95 1.38 2.395 ;
      RECT 1.475 0.425 1.805 0.965 ;
      RECT 0.115 1.11 1.305 1.28 ;
      RECT 0.115 0.35 0.365 1.11 ;
      RECT 1.055 0.35 1.305 1.11 ;
      RECT 1.615 1.975 2.565 2.225 ;
      RECT 1.615 1.135 2.375 1.305 ;
      RECT 2.045 0.595 2.375 1.135 ;
      RECT 1.615 1.78 1.785 1.975 ;
      RECT 1.455 1.45 1.785 1.78 ;
      RECT 1.615 1.305 1.785 1.45 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 3.955 1.82 4.205 3.245 ;
      RECT 1.585 2.735 1.94 3.245 ;
      RECT 2.77 2.735 3.22 3.245 ;
      RECT 0.12 1.95 0.45 3.245 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 3.94 0.085 4.19 1.13 ;
      RECT 0.545 0.085 0.875 0.94 ;
      RECT 2.885 0.085 3.215 0.965 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o2bb2a_2

MACRO scs8ls_o2bb2a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.415 1.35 4.745 1.78 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END A1N

  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.845 1.35 4.195 1.78 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END A2N

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.26 1.115 1.77 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.47 1.45 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B2

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.255 0.81 6.585 1.05 ;
        RECT 6.255 1.05 6.585 1.72 ;
        RECT 5.255 0.35 5.585 0.81 ;
        RECT 6.255 0.35 6.585 0.81 ;
        RECT 5.255 1.72 6.585 1.89 ;
        RECT 5.255 1.89 5.585 2.98 ;
        RECT 6.255 1.89 6.585 2.98 ;
    END
    ANTENNADIFFAREA 1.3113 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.085 2.905 2.315 3.075 ;
      RECT 1.985 2.29 2.315 2.905 ;
      RECT 1.085 2.12 1.415 2.905 ;
      RECT 0.185 1.95 1.415 2.12 ;
      RECT 0.185 2.12 0.515 2.98 ;
      RECT 0.185 1.94 0.515 1.95 ;
      RECT 0.115 0.92 3.335 1.09 ;
      RECT 1.115 0.78 3.335 0.92 ;
      RECT 0.115 0.35 0.445 0.92 ;
      RECT 3.005 0.595 3.335 0.78 ;
      RECT 1.115 0.35 1.445 0.78 ;
      RECT 3.505 1.95 4.465 2.28 ;
      RECT 3.505 0.96 4.03 1.13 ;
      RECT 3.7 0.635 4.03 0.96 ;
      RECT 3.505 1.63 3.675 1.95 ;
      RECT 2.49 1.3 3.675 1.63 ;
      RECT 3.505 1.13 3.675 1.3 ;
      RECT 4.915 1.22 6.065 1.55 ;
      RECT 3.165 2.45 5.085 2.62 ;
      RECT 4.915 1.55 5.085 2.45 ;
      RECT 4.915 1.12 5.085 1.22 ;
      RECT 4.2 0.95 5.085 1.12 ;
      RECT 4.2 0.425 4.37 0.95 ;
      RECT 2.505 0.255 4.37 0.425 ;
      RECT 3.165 2.15 3.335 2.45 ;
      RECT 2.995 2.12 3.335 2.15 ;
      RECT 1.615 1.95 3.335 2.12 ;
      RECT 1.615 2.12 1.785 2.735 ;
      RECT 2.995 1.82 3.335 1.95 ;
      RECT 2.505 0.425 2.835 0.61 ;
      RECT 0 -0.085 7.2 0.085 ;
      RECT 6.755 0.085 7.085 1.13 ;
      RECT 0.615 0.085 0.945 0.75 ;
      RECT 1.615 0.085 1.945 0.61 ;
      RECT 4.54 0.085 5.08 0.78 ;
      RECT 5.755 0.085 6.085 0.64 ;
      RECT 0 3.245 7.2 3.415 ;
      RECT 6.755 1.82 7.085 3.245 ;
      RECT 3.6 2.79 3.93 3.245 ;
      RECT 4.67 2.79 5 3.245 ;
      RECT 2.545 2.32 2.875 3.245 ;
      RECT 0.715 2.29 0.885 3.245 ;
      RECT 5.755 2.06 6.085 3.245 ;
    LAYER mcon ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_o2bb2a_4

MACRO scs8ls_o2bb2ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.12 1.1 1.45 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END A2N

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.3 3.255 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.435 1.51 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END A1N

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.225 1.3 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.86 1.95 2.315 2.98 ;
        RECT 1.86 1.18 2.03 1.95 ;
        RECT 1.61 1.01 2.03 1.18 ;
        RECT 1.61 0.35 1.86 1.01 ;
    END
    ANTENNADIFFAREA 0.5469 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.64 1.62 1.69 1.79 ;
      RECT 1.27 1.35 1.69 1.62 ;
      RECT 0.64 1.79 0.97 2.775 ;
      RECT 1.27 0.95 1.44 1.35 ;
      RECT 0.935 0.35 1.44 0.95 ;
      RECT 2.2 0.96 3.22 1.13 ;
      RECT 2.2 0.84 2.37 0.96 ;
      RECT 2.89 0.35 3.22 0.96 ;
      RECT 2.03 0.445 2.37 0.84 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.54 0.085 2.71 0.79 ;
      RECT 0.115 0.085 0.445 0.95 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.995 1.95 3.245 3.245 ;
      RECT 1.14 1.975 1.69 3.245 ;
      RECT 0.14 1.895 0.47 3.245 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_o2bb2ai_1

MACRO scs8ls_o2bb2ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.63 0.355 2.415 ;
        RECT 0.125 1.3 0.48 1.63 ;
        RECT 0.125 2.415 0.82 2.45 ;
        RECT 0.125 2.45 2.335 2.585 ;
        RECT 0.65 2.585 2.335 2.62 ;
        RECT 2.165 1.68 2.335 2.45 ;
        RECT 1.965 1.35 2.335 1.68 ;
    END
    ANTENNAGATEAREA 0.444 ;
  END A1N

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.35 5.495 1.72 ;
        RECT 3.695 1.72 5.495 1.78 ;
        RECT 3.695 1.78 5.095 1.89 ;
        RECT 3.695 1.35 4.025 1.72 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3 0.595 3.29 1.13 ;
        RECT 3.005 1.13 3.29 2.06 ;
        RECT 3.005 2.06 4.695 2.23 ;
        RECT 3.005 2.23 3.29 2.98 ;
        RECT 4.465 2.23 4.695 2.735 ;
    END
    ANTENNADIFFAREA 0.896 ;
  END Y

  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.375 1.445 1.795 1.78 ;
    END
    ANTENNAGATEAREA 0.444 ;
  END A2N

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.345 1.18 4.675 1.55 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.65 1.105 2.675 1.18 ;
      RECT 2.505 1.18 2.675 1.3 ;
      RECT 1.155 1.01 2.675 1.105 ;
      RECT 2.505 1.3 2.835 1.63 ;
      RECT 0.65 1.18 1.405 1.275 ;
      RECT 1.155 0.605 1.405 1.01 ;
      RECT 1.72 2.245 1.995 2.28 ;
      RECT 0.65 1.95 1.995 2.245 ;
      RECT 0.65 1.275 0.98 1.95 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 3.96 0.085 4.29 0.67 ;
      RECT 4.87 0.085 5.215 0.6 ;
      RECT 0.145 0.085 0.475 1.03 ;
      RECT 2.08 0.085 2.34 0.825 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 5.395 1.95 5.645 3.245 ;
      RECT 2.505 1.82 2.835 3.245 ;
      RECT 0.115 2.755 0.445 3.245 ;
      RECT 1.185 2.79 1.515 3.245 ;
      RECT 3.46 2.4 3.79 3.245 ;
      RECT 3.965 2.905 5.195 3.075 ;
      RECT 4.865 2.06 5.195 2.905 ;
      RECT 3.965 2.4 4.295 2.905 ;
      RECT 0.645 0.425 0.975 0.935 ;
      RECT 0.645 0.255 1.91 0.425 ;
      RECT 1.58 0.425 1.91 0.825 ;
      RECT 3.46 1.01 3.79 1.13 ;
      RECT 3.46 0.84 5.645 1.01 ;
      RECT 5.315 1.01 5.645 1.13 ;
      RECT 3.46 0.425 3.79 0.84 ;
      RECT 4.47 0.77 5.645 0.84 ;
      RECT 2.57 0.255 3.79 0.425 ;
      RECT 4.47 0.35 4.69 0.77 ;
      RECT 5.395 0.35 5.645 0.77 ;
      RECT 2.57 0.425 2.82 0.825 ;
    LAYER mcon ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_o2bb2ai_2

MACRO scs8ls_o2bb2ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.35 7.64 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.15 1.35 9.955 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B1

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.935 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1N

  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.225 1.35 3.235 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2N

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.055 1.97 7.725 2.12 ;
        RECT 5.055 2.12 5.635 2.15 ;
        RECT 6.495 2.12 6.825 2.735 ;
        RECT 7.395 2.12 7.725 2.735 ;
        RECT 4.155 1.95 7.725 1.97 ;
        RECT 4.155 1.8 5.715 1.95 ;
        RECT 5.055 2.15 5.305 2.98 ;
        RECT 4.155 1.97 4.485 2.98 ;
        RECT 5.545 1.13 5.715 1.8 ;
        RECT 4.695 0.96 5.885 1.13 ;
        RECT 4.695 0.595 5.025 0.96 ;
        RECT 5.545 0.595 5.885 0.96 ;
    END
    ANTENNADIFFAREA 1.7584 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.115 1.01 2.095 1.18 ;
      RECT 1.925 0.425 2.095 1.01 ;
      RECT 0.115 0.35 0.365 1.01 ;
      RECT 1.055 0.35 1.235 1.01 ;
      RECT 1.925 0.255 4.035 0.425 ;
      RECT 2.775 0.425 3.105 0.84 ;
      RECT 3.785 0.425 4.035 1.13 ;
      RECT 6.065 1.01 9.965 1.18 ;
      RECT 6.065 0.425 6.235 1.01 ;
      RECT 6.915 0.35 7.165 1.01 ;
      RECT 7.845 0.35 8.095 1.01 ;
      RECT 8.785 0.35 9.035 1.01 ;
      RECT 9.715 0.35 9.965 1.01 ;
      RECT 4.265 0.255 6.235 0.425 ;
      RECT 4.265 0.425 4.515 1.13 ;
      RECT 5.205 0.425 5.375 0.79 ;
      RECT 3.415 1.3 5.375 1.63 ;
      RECT 0.555 1.95 3.585 2.12 ;
      RECT 2.355 2.12 2.685 2.98 ;
      RECT 3.255 2.12 3.585 2.98 ;
      RECT 3.415 1.63 3.585 1.95 ;
      RECT 3.415 1.18 3.605 1.3 ;
      RECT 2.275 1.01 3.605 1.18 ;
      RECT 2.275 0.595 2.605 1.01 ;
      RECT 3.275 0.595 3.605 1.01 ;
      RECT 0.555 2.12 0.885 2.98 ;
      RECT 1.455 2.12 1.785 2.98 ;
      RECT 6.045 2.905 8.11 3.075 ;
      RECT 7.91 2.12 8.11 2.905 ;
      RECT 7.91 1.95 9.975 2.12 ;
      RECT 8.745 2.12 9.075 2.98 ;
      RECT 9.645 2.12 9.975 2.98 ;
      RECT 6.045 2.29 6.31 2.905 ;
      RECT 7.01 2.29 7.21 2.905 ;
      RECT 0 3.245 10.08 3.415 ;
      RECT 8.295 2.29 8.56 3.245 ;
      RECT 9.26 2.29 9.465 3.245 ;
      RECT 1.085 2.29 1.255 3.245 ;
      RECT 1.985 2.29 2.155 3.245 ;
      RECT 2.885 2.29 3.055 3.245 ;
      RECT 0.105 1.95 0.355 3.245 ;
      RECT 3.785 1.82 3.955 3.245 ;
      RECT 4.685 2.14 4.855 3.245 ;
      RECT 5.505 2.32 5.835 3.245 ;
      RECT 0 -0.085 10.08 0.085 ;
      RECT 6.415 0.085 6.745 0.83 ;
      RECT 7.345 0.085 7.675 0.83 ;
      RECT 8.275 0.085 8.605 0.83 ;
      RECT 9.205 0.085 9.535 0.83 ;
      RECT 0.545 0.085 0.875 0.84 ;
      RECT 1.415 0.085 1.745 0.84 ;
    LAYER mcon ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
  END
END scs8ls_o2bb2ai_4

MACRO scs8ls_o311a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.87 0.35 4.235 1.13 ;
        RECT 4.065 1.13 4.235 1.96 ;
        RECT 3.855 1.96 4.235 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.015 1.12 3.385 1.45 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455 1.14 1.805 1.47 ;
        RECT 1.635 1.47 1.805 2.32 ;
        RECT 1.635 2.32 2.845 2.49 ;
        RECT 2.515 1.445 2.845 2.32 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975 1.12 2.305 2.15 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.92 1.14 1.285 1.47 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.14 0.41 1.47 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END C1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.06 0.61 1.39 0.97 ;
      RECT 1.06 0.28 3.18 0.61 ;
      RECT 3.015 1.62 3.895 1.79 ;
      RECT 3.595 1.35 3.895 1.62 ;
      RECT 1.135 2.785 3.185 2.955 ;
      RECT 3.015 1.79 3.185 2.785 ;
      RECT 0.135 1.64 1.465 1.81 ;
      RECT 1.135 1.81 1.465 2.785 ;
      RECT 0.135 1.81 0.465 2.955 ;
      RECT 0.58 0.97 0.75 1.64 ;
      RECT 0.2 0.8 0.75 0.97 ;
      RECT 0.2 0.35 0.53 0.8 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 1.56 0.78 3.69 0.95 ;
      RECT 3.36 0.085 3.69 0.78 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 3.355 1.96 3.685 3.245 ;
      RECT 0.635 1.98 0.965 3.245 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_o311a_1

MACRO scs8ls_o311a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.435 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END C1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 1.35 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.35 1.815 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025 1.35 2.355 2.89 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.35 2.925 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.435 0.81 4.195 1.05 ;
        RECT 3.965 1.05 4.195 1.72 ;
        RECT 3.435 0.35 3.685 0.81 ;
        RECT 3.33 1.72 4.195 1.89 ;
        RECT 3.33 1.89 3.66 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.18 0.67 2.66 0.84 ;
      RECT 1.18 0.35 1.51 0.67 ;
      RECT 2.33 0.35 2.66 0.67 ;
      RECT 3.095 1.22 3.51 1.55 ;
      RECT 0.605 1.01 3.265 1.18 ;
      RECT 3.095 1.18 3.265 1.22 ;
      RECT 0.225 1.95 1.665 2.12 ;
      RECT 1.335 2.12 1.665 2.98 ;
      RECT 0.225 2.12 0.605 2.86 ;
      RECT 0.225 1.82 0.775 1.95 ;
      RECT 0.605 1.18 0.775 1.82 ;
      RECT 0.205 0.35 0.775 1.01 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 3.83 2.06 4.16 3.245 ;
      RECT 2.745 1.95 3.075 3.245 ;
      RECT 0.775 2.29 1.105 3.245 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 3.855 0.085 4.205 0.6 ;
      RECT 1.69 0.085 2.15 0.5 ;
      RECT 2.83 0.085 3.16 0.84 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o311a_2

MACRO scs8ls_o311a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.14 0.945 1.31 ;
        RECT 0.125 1.31 0.355 1.48 ;
        RECT 0.615 1.05 0.945 1.14 ;
        RECT 0.125 1.48 0.895 1.65 ;
        RECT 0.615 0.88 2.07 1.05 ;
        RECT 0.565 1.65 0.895 1.72 ;
        RECT 0.615 0.35 0.945 0.88 ;
        RECT 1.74 0.35 2.07 0.88 ;
        RECT 0.565 1.72 1.895 1.89 ;
        RECT 0.565 1.89 0.895 2.98 ;
        RECT 1.565 1.89 1.895 2.98 ;
    END
    ANTENNADIFFAREA 1.3454 ;
  END X

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.105 1.47 8.035 1.8 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.525 1.22 8.535 1.3 ;
        RECT 8.205 1.3 8.535 1.78 ;
        RECT 6.525 1.3 6.935 1.55 ;
        RECT 6.765 1.13 8.535 1.22 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.87 1.42 6.2 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.64 5.36 1.8 ;
        RECT 3.995 1.47 5.36 1.64 ;
        RECT 3.995 1.265 4.165 1.47 ;
        RECT 2.505 1.22 4.165 1.265 ;
        RECT 2.505 1.265 2.91 1.55 ;
        RECT 2.74 1.095 4.165 1.22 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.435 3.825 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END C1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 6.22 2.96 8.525 3.075 ;
      RECT 5.15 2.905 8.525 2.96 ;
      RECT 5.15 2.71 6.55 2.905 ;
      RECT 8.195 1.97 8.525 2.905 ;
      RECT 6.265 0.96 6.595 1.05 ;
      RECT 5.265 0.79 8.525 0.96 ;
      RECT 5.265 0.425 5.595 0.79 ;
      RECT 6.265 0.37 6.595 0.79 ;
      RECT 7.265 0.35 7.595 0.79 ;
      RECT 8.275 0.35 8.525 0.79 ;
      RECT 2.8 0.255 5.595 0.425 ;
      RECT 2.8 0.425 3.13 0.925 ;
      RECT 3.3 0.765 4.075 0.925 ;
      RECT 3.3 0.595 5.095 0.765 ;
      RECT 4.765 0.765 5.095 0.96 ;
      RECT 6.72 2.565 8.025 2.735 ;
      RECT 7.775 1.97 8.025 2.565 ;
      RECT 4.09 2.12 6.1 2.14 ;
      RECT 5.75 2.14 6.1 2.2 ;
      RECT 2.655 1.97 6.1 2.12 ;
      RECT 5.53 1.95 6.1 1.97 ;
      RECT 5.53 1.3 5.7 1.95 ;
      RECT 4.335 1.13 5.7 1.3 ;
      RECT 4.09 2.14 4.42 2.98 ;
      RECT 2.655 1.95 4.42 1.97 ;
      RECT 4.09 1.94 4.42 1.95 ;
      RECT 4.335 0.935 4.585 1.13 ;
      RECT 2.095 1.55 2.265 1.72 ;
      RECT 1.255 1.22 2.265 1.55 ;
      RECT 2.655 2.12 2.985 2.98 ;
      RECT 2.655 1.89 2.985 1.95 ;
      RECT 2.095 1.72 2.985 1.89 ;
      RECT 0 -0.085 8.64 0.085 ;
      RECT 2.24 0.085 2.57 1.05 ;
      RECT 5.765 0.085 6.095 0.62 ;
      RECT 6.765 0.085 7.095 0.62 ;
      RECT 7.765 0.085 8.095 0.62 ;
      RECT 0.115 0.085 0.445 0.97 ;
      RECT 1.115 0.085 1.57 0.68 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 4.59 2.54 4.92 3.245 ;
      RECT 3.225 2.29 3.92 3.245 ;
      RECT 2.15 2.06 2.48 3.245 ;
      RECT 4.59 2.395 6.55 2.54 ;
      RECT 4.59 2.37 7.575 2.395 ;
      RECT 4.59 2.31 4.92 2.37 ;
      RECT 6.38 1.97 7.575 2.37 ;
      RECT 0.115 1.82 0.365 3.245 ;
      RECT 1.065 2.06 1.395 3.245 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
  END
END scs8ls_o311a_4

MACRO scs8ls_o311ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515 1.18 1.845 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A3

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.805 1.89 3.235 2.98 ;
        RECT 1.785 1.72 3.235 1.89 ;
        RECT 1.785 1.89 2.115 2.98 ;
        RECT 2.585 1.01 2.755 1.72 ;
        RECT 2.585 0.35 3.11 1.01 ;
    END
    ANTENNADIFFAREA 1.0117 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.18 2.415 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.18 3.255 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END C1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 0.705 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 1.35 1.315 2.89 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.615 1.01 0.945 1.13 ;
      RECT 0.615 0.84 2.22 1.01 ;
      RECT 0.615 0.35 0.945 0.84 ;
      RECT 1.89 0.33 2.22 0.84 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.285 2.06 2.615 3.245 ;
      RECT 0.225 1.95 0.555 3.245 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 0.115 0.085 0.445 1.13 ;
      RECT 1.115 0.085 1.675 0.65 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o311ai_1

MACRO scs8ls_o311ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.4 0.595 4.705 0.96 ;
        RECT 4.4 0.96 5.645 1.13 ;
        RECT 4.4 1.13 4.73 1.95 ;
        RECT 5.395 0.35 5.645 0.96 ;
        RECT 2.6 1.95 5.63 2.12 ;
        RECT 2.6 2.12 2.93 2.735 ;
        RECT 3.5 2.12 3.75 2.98 ;
        RECT 4.48 2.12 4.65 2.98 ;
        RECT 5.3 2.12 5.63 2.98 ;
    END
    ANTENNADIFFAREA 1.7546 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.35 4.195 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.3 5.635 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END C1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.35 3.235 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.35 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.395 0.255 5.215 0.425 ;
      RECT 4.885 0.425 5.215 0.79 ;
      RECT 3.395 0.425 3.725 0.84 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 0.65 2.29 0.9 3.245 ;
      RECT 3.95 2.29 4.28 3.245 ;
      RECT 4.85 2.29 5.1 3.245 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 0.545 0.085 0.875 0.84 ;
      RECT 1.535 0.085 1.865 0.84 ;
      RECT 2.465 0.085 2.795 0.84 ;
      RECT 0.12 2.12 0.45 2.98 ;
      RECT 0.12 1.95 2.37 2.12 ;
      RECT 1.07 2.12 1.4 2.98 ;
      RECT 2.12 2.12 2.37 2.735 ;
      RECT 1.59 2.905 3.3 3.075 ;
      RECT 3.13 2.29 3.3 2.905 ;
      RECT 1.59 2.29 1.92 2.905 ;
      RECT 0.115 1.01 4.225 1.18 ;
      RECT 3.895 0.595 4.225 1.01 ;
      RECT 0.115 0.35 0.365 1.01 ;
      RECT 1.115 0.35 1.365 1.01 ;
      RECT 2.045 0.35 2.295 1.01 ;
      RECT 2.975 0.35 3.225 1.01 ;
    LAYER mcon ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o311ai_2

MACRO scs8ls_o311ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 11.04 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.165 1.35 10.435 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.765 1.35 7.775 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.185 1.64 6.195 1.78 ;
        RECT 4.485 1.43 6.195 1.64 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.245 1.43 4.195 1.78 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.3 1.24 1.78 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END C1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.26 6.595 1.95 ;
        RECT 0.74 1.95 6.595 2.12 ;
        RECT 1.41 1.1 6.595 1.26 ;
        RECT 0.74 2.12 1.07 2.98 ;
        RECT 1.74 2.12 2.07 2.98 ;
        RECT 4.685 2.12 5.015 2.735 ;
        RECT 5.685 2.12 6.015 2.735 ;
        RECT 1.74 1.82 2.07 1.95 ;
        RECT 4.685 1.82 5.015 1.95 ;
        RECT 0.545 1.09 6.595 1.1 ;
        RECT 0.545 0.77 1.74 1.09 ;
    END
    ANTENNADIFFAREA 2.2717 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.04 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.04 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 8.725 0.96 10.415 1.13 ;
      RECT 10.165 0.35 10.415 0.96 ;
      RECT 7.945 1.3 8.975 1.47 ;
      RECT 7.945 1.18 8.115 1.3 ;
      RECT 8.725 1.13 8.975 1.3 ;
      RECT 6.89 1.01 8.115 1.18 ;
      RECT 6.89 0.92 7.14 1.01 ;
      RECT 7.945 0.35 8.115 1.01 ;
      RECT 8.725 0.35 8.975 0.96 ;
      RECT 4.07 0.75 7.14 0.92 ;
      RECT 6.89 0.35 7.14 0.75 ;
      RECT 4.92 0.35 5.17 0.75 ;
      RECT 5.86 0.35 6.19 0.75 ;
      RECT 4.07 0.58 4.24 0.75 ;
      RECT 2.27 0.33 4.24 0.58 ;
      RECT 1.92 0.75 3.9 0.92 ;
      RECT 1.92 0.6 2.09 0.75 ;
      RECT 0.115 0.35 2.09 0.6 ;
      RECT 0.115 0.6 0.365 1.13 ;
      RECT 7.785 2.15 8.065 2.735 ;
      RECT 7.785 2.12 10.475 2.15 ;
      RECT 9.295 2.15 9.525 2.98 ;
      RECT 10.195 2.15 10.475 2.98 ;
      RECT 6.785 1.95 10.475 2.12 ;
      RECT 6.785 2.12 7.115 2.735 ;
      RECT 4.185 2.905 8.565 3.075 ;
      RECT 8.235 2.33 8.565 2.905 ;
      RECT 6.285 2.29 6.615 2.905 ;
      RECT 7.285 2.29 7.615 2.905 ;
      RECT 4.185 2.29 4.515 2.905 ;
      RECT 5.185 2.29 5.515 2.905 ;
      RECT 4.41 0.085 4.74 0.58 ;
      RECT 0 -0.085 11.04 0.085 ;
      RECT 5.35 0.085 5.68 0.58 ;
      RECT 6.37 0.085 6.71 0.58 ;
      RECT 7.32 0.085 7.65 0.825 ;
      RECT 8.295 0.085 8.545 1.13 ;
      RECT 9.155 0.085 9.995 0.79 ;
      RECT 10.595 0.085 10.925 1.13 ;
      RECT 0 3.245 11.04 3.415 ;
      RECT 8.795 2.33 9.125 3.245 ;
      RECT 9.695 2.33 10.025 3.245 ;
      RECT 10.675 1.82 10.925 3.245 ;
      RECT 0.115 1.95 0.445 3.245 ;
      RECT 1.24 2.29 1.57 3.245 ;
      RECT 2.24 2.29 3.905 3.245 ;
    LAYER mcon ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
  END
END scs8ls_o311ai_4

MACRO scs8ls_o31a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.82 0.455 2.98 ;
        RECT 0.085 1.13 0.255 1.82 ;
        RECT 0.085 0.35 0.445 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 2.375 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A3

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.35 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.3 1.835 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.545 1.35 2.915 1.78 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END B1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.125 0.96 2.745 1.13 ;
      RECT 1.125 0.45 1.46 0.96 ;
      RECT 2.415 0.45 2.745 0.96 ;
      RECT 0.625 1.95 3.255 2.12 ;
      RECT 3.085 1.13 3.255 1.95 ;
      RECT 2.915 0.45 3.255 1.13 ;
      RECT 2.195 2.12 2.525 2.88 ;
      RECT 0.625 1.65 0.795 1.95 ;
      RECT 0.425 1.32 0.795 1.65 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 0.625 2.29 1.09 3.245 ;
      RECT 2.735 2.29 3.05 3.245 ;
      RECT 0.615 0.085 0.945 1.13 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 1.765 0.085 2.13 0.78 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o31a_1

MACRO scs8ls_o31a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.82 0.95 2.15 ;
        RECT 0.775 1.13 0.945 1.82 ;
        RECT 0.615 0.35 0.945 1.13 ;
    END
    ANTENNADIFFAREA 0.6048 ;
  END X

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415 1.35 1.795 2.15 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 1.47 2.315 2.15 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.18 2.885 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395 1.3 3.725 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.615 0.94 1.945 1.13 ;
      RECT 1.615 0.79 2.85 0.94 ;
      RECT 1.615 0.77 3.225 0.79 ;
      RECT 2.68 0.46 3.225 0.77 ;
      RECT 1.615 0.35 1.945 0.77 ;
      RECT 3.055 0.96 3.725 1.13 ;
      RECT 3.395 0.35 3.725 0.96 ;
      RECT 2.765 2.49 3.225 2.98 ;
      RECT 0.225 2.32 3.225 2.49 ;
      RECT 2.765 1.94 3.225 2.32 ;
      RECT 3.055 1.13 3.225 1.94 ;
      RECT 0.225 1.65 0.395 2.32 ;
      RECT 0.225 1.32 0.605 1.65 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 1.115 0.085 1.445 1.13 ;
      RECT 2.115 0.085 2.51 0.6 ;
      RECT 0.115 0.085 0.445 1.13 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 3.395 1.95 3.725 3.245 ;
      RECT 1.07 2.66 1.595 3.245 ;
      RECT 0.115 2.66 0.445 3.245 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_o31a_2

MACRO scs8ls_o31a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575 0.35 0.905 0.96 ;
        RECT 0.575 0.96 1.7 1.13 ;
        RECT 0.575 1.13 0.835 1.8 ;
        RECT 1.45 0.35 1.7 0.96 ;
        RECT 0.575 1.8 1.81 1.97 ;
        RECT 0.575 1.97 0.835 2.98 ;
        RECT 1.48 1.97 1.81 2.98 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END X

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.47 3.235 2.15 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.455 5.155 1.785 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A3

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405 1.455 5.875 1.785 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.115 1.455 6.595 1.785 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.45 1.115 6.58 1.285 ;
      RECT 4.39 0.605 4.64 1.115 ;
      RECT 5.32 0.605 5.57 1.115 ;
      RECT 6.25 0.605 6.58 1.115 ;
      RECT 3.45 0.435 3.78 1.115 ;
      RECT 2.44 0.265 3.78 0.435 ;
      RECT 2.44 0.435 2.77 0.96 ;
      RECT 4.825 2.465 5.075 2.98 ;
      RECT 4.825 2.295 6.105 2.465 ;
      RECT 5.775 2.465 6.105 2.98 ;
      RECT 2.465 2.375 4.255 2.545 ;
      RECT 3.925 2.545 4.255 2.98 ;
      RECT 2.545 1.13 3.27 1.3 ;
      RECT 2.94 0.605 3.27 1.13 ;
      RECT 2.465 2.545 2.715 2.98 ;
      RECT 2.465 1.63 2.715 2.375 ;
      RECT 1.005 1.3 2.715 1.63 ;
      RECT 4.435 2.205 4.645 2.98 ;
      RECT 3.475 2.125 4.645 2.205 ;
      RECT 3.475 1.955 6.605 2.125 ;
      RECT 6.275 2.125 6.605 2.98 ;
      RECT 0 3.245 6.72 3.415 ;
      RECT 2.915 2.715 3.245 3.245 ;
      RECT 5.275 2.635 5.605 3.245 ;
      RECT 2.01 1.82 2.26 3.245 ;
      RECT 0.13 1.82 0.38 3.245 ;
      RECT 1.03 2.14 1.28 3.245 ;
      RECT 0 -0.085 6.72 0.085 ;
      RECT 1.88 0.085 2.21 1.13 ;
      RECT 3.96 0.085 4.21 0.945 ;
      RECT 4.82 0.085 5.15 0.945 ;
      RECT 5.75 0.085 6.08 0.945 ;
      RECT 0.145 0.085 0.395 1.13 ;
      RECT 1.085 0.085 1.255 0.79 ;
    LAYER mcon ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
  END
END scs8ls_o31a_4

MACRO scs8ls_o31ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.35 1.95 2.23 2.98 ;
        RECT 1.35 1.13 1.52 1.95 ;
        RECT 1.35 0.96 2.765 1.13 ;
        RECT 2.435 0.35 2.765 0.96 ;
    END
    ANTENNADIFFAREA 1.0207 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.435 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.3 2.775 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.3 1.18 2.89 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.69 1.35 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A3

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.625 0.62 2.265 0.79 ;
      RECT 1.935 0.35 2.265 0.62 ;
      RECT 0.625 0.79 0.875 1.13 ;
      RECT 0.625 0.35 0.875 0.62 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 2.41 1.95 2.74 3.245 ;
      RECT 0.13 1.82 0.38 3.245 ;
      RECT 0 -0.085 2.88 0.085 ;
      RECT 0.115 0.085 0.445 1.01 ;
      RECT 1.055 0.085 1.755 0.45 ;
    LAYER mcon ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o31ai_1

MACRO scs8ls_o31ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.455 2.12 3.785 2.98 ;
        RECT 2.505 2.02 3.785 2.12 ;
        RECT 2.505 2.12 2.755 2.735 ;
        RECT 2.505 1.95 4.685 2.02 ;
        RECT 4.355 2.02 4.685 2.98 ;
        RECT 3.615 1.85 4.685 1.95 ;
        RECT 2.505 1.82 2.835 1.95 ;
        RECT 2.665 1.18 2.835 1.82 ;
        RECT 2.665 1.01 4.18 1.18 ;
        RECT 3.85 0.61 4.18 1.01 ;
    END
    ANTENNADIFFAREA 1.297 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.35 3.445 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.365 1.18 4.695 1.35 ;
        RECT 3.685 1.35 4.695 1.68 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.35 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.55 2.905 3.285 3.075 ;
      RECT 2.955 2.29 3.285 2.905 ;
      RECT 1.55 2.29 1.72 2.905 ;
      RECT 3.42 0.255 4.68 0.425 ;
      RECT 4.35 0.425 4.68 1.01 ;
      RECT 0.115 1.01 2.445 1.18 ;
      RECT 2.115 0.84 2.445 1.01 ;
      RECT 0.115 0.35 0.445 1.01 ;
      RECT 1.115 0.35 1.445 1.01 ;
      RECT 2.115 0.35 2.445 0.67 ;
      RECT 2.115 0.67 3.67 0.84 ;
      RECT 3.42 0.425 3.67 0.67 ;
      RECT 0.12 2.12 0.37 2.98 ;
      RECT 0.12 1.95 2.25 2.12 ;
      RECT 1.02 2.12 1.35 2.98 ;
      RECT 1.92 2.12 2.25 2.735 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 0.57 2.29 0.82 3.245 ;
      RECT 3.985 2.19 4.155 3.245 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 0.615 0.085 0.945 0.825 ;
      RECT 1.615 0.085 1.945 0.825 ;
      RECT 2.625 0.085 3.24 0.5 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o31ai_2

MACRO scs8ls_o31ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.795 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.35 3.715 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.835 1.35 6.115 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.35 7.79 1.78 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.55 4.665 1.95 ;
        RECT 3.965 1.95 8.525 2.12 ;
        RECT 4.495 1.18 4.665 1.55 ;
        RECT 3.965 2.12 4.97 2.15 ;
        RECT 5.6 2.12 5.93 2.735 ;
        RECT 6.55 2.12 6.88 2.98 ;
        RECT 8.195 2.12 8.525 2.98 ;
        RECT 8.195 1.82 8.525 1.95 ;
        RECT 4.495 1.01 8.095 1.18 ;
        RECT 4.7 2.15 4.97 2.735 ;
        RECT 6.905 0.92 8.095 1.01 ;
    END
    ANTENNADIFFAREA 1.8032 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 6.475 0.39 8.525 0.56 ;
      RECT 7.335 0.56 7.665 0.75 ;
      RECT 8.265 0.56 8.525 1.17 ;
      RECT 0.115 1.01 4.325 1.18 ;
      RECT 0.115 0.92 2.305 1.01 ;
      RECT 4.155 0.84 4.325 1.01 ;
      RECT 3.145 0.39 3.475 1.01 ;
      RECT 0.115 0.39 0.445 0.92 ;
      RECT 1.975 0.39 2.305 0.92 ;
      RECT 4.155 0.39 4.325 0.67 ;
      RECT 4.155 0.75 5.775 0.84 ;
      RECT 4.155 0.67 6.805 0.75 ;
      RECT 5.445 0.58 6.805 0.67 ;
      RECT 6.475 0.56 6.805 0.58 ;
      RECT 5.445 0.39 5.775 0.58 ;
      RECT 2.97 2.37 4.47 2.54 ;
      RECT 4.14 2.54 4.47 2.735 ;
      RECT 2.97 2.54 3.3 2.735 ;
      RECT 2.97 2.12 3.3 2.37 ;
      RECT 0.12 1.95 3.3 2.12 ;
      RECT 0.12 2.12 0.37 2.98 ;
      RECT 1.1 2.12 1.27 2.98 ;
      RECT 1.97 2.12 2.3 2.98 ;
      RECT 1.97 1.82 2.3 1.95 ;
      RECT 2.47 2.905 6.38 3.075 ;
      RECT 6.13 2.29 6.38 2.905 ;
      RECT 3.64 2.71 3.97 2.905 ;
      RECT 2.47 2.29 2.8 2.905 ;
      RECT 5.15 2.29 5.4 2.905 ;
      RECT 0.615 0.085 0.945 0.75 ;
      RECT 0 -0.085 8.64 0.085 ;
      RECT 1.475 0.085 1.805 0.75 ;
      RECT 2.495 0.085 2.96 0.805 ;
      RECT 3.645 0.085 3.975 0.84 ;
      RECT 4.585 0.085 5.265 0.5 ;
      RECT 5.955 0.085 6.295 0.41 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 0.57 2.29 0.9 3.245 ;
      RECT 1.47 2.29 1.8 3.245 ;
      RECT 7.05 2.29 8.025 3.245 ;
    LAYER mcon ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
  END
END scs8ls_o31ai_4

MACRO scs8ls_o32a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.35 0.56 1.13 ;
        RECT 0.085 1.13 0.255 1.82 ;
        RECT 0.085 1.82 0.445 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.535 1.35 2.895 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.035 1.35 2.365 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495 1.35 1.825 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955 1.35 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.41 1.18 3.735 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.23 1.01 2.56 1.18 ;
      RECT 2.23 0.52 2.56 1.01 ;
      RECT 1.23 0.35 1.56 1.01 ;
      RECT 2.23 0.34 3.655 0.52 ;
      RECT 3.405 0.52 3.655 1.01 ;
      RECT 2.205 2.12 2.595 2.88 ;
      RECT 0.615 1.95 3.235 2.12 ;
      RECT 3.065 1.18 3.235 1.95 ;
      RECT 2.73 1.01 3.235 1.18 ;
      RECT 2.73 0.7 3.225 1.01 ;
      RECT 0.615 1.65 0.785 1.95 ;
      RECT 0.425 1.32 0.785 1.65 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 0.615 2.29 0.945 3.245 ;
      RECT 3.32 2.29 3.65 3.245 ;
      RECT 3.41 1.97 3.65 2.29 ;
      RECT 0.73 0.085 1.06 1.03 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 1.73 0.085 2.06 0.82 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o32a_1

MACRO scs8ls_o32a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 1.82 0.895 2.98 ;
        RECT 0.535 1.13 0.705 1.82 ;
        RECT 0.535 0.96 1.05 1.13 ;
        RECT 0.72 0.35 1.05 0.96 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.095 1.35 3.715 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.355 1.18 4.685 2.89 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.35 2.855 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 1.35 2.315 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415 1.35 1.795 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.72 1.01 3.05 1.18 ;
      RECT 2.72 0.52 3.05 1.01 ;
      RECT 1.72 0.35 2.05 1.01 ;
      RECT 2.72 0.35 4.615 0.52 ;
      RECT 4.355 0.52 4.615 1.01 ;
      RECT 2.675 2.12 3.11 2.88 ;
      RECT 1.065 1.95 4.185 2.12 ;
      RECT 4.015 1.045 4.185 1.95 ;
      RECT 3.22 0.715 4.185 1.045 ;
      RECT 1.065 1.65 1.235 1.95 ;
      RECT 0.875 1.32 1.235 1.65 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 1.065 2.29 1.6 3.245 ;
      RECT 3.815 2.29 4.145 3.245 ;
      RECT 0.115 1.82 0.365 3.245 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 1.22 0.085 1.55 1.13 ;
      RECT 2.22 0.085 2.55 0.84 ;
      RECT 0.115 0.79 0.365 1.14 ;
      RECT 0.115 0.085 0.54 0.79 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o32a_2

MACRO scs8ls_o32a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.45 2.855 1.78 ;
        RECT 2.685 1.78 2.855 2.36 ;
        RECT 2.685 2.36 5.905 2.53 ;
        RECT 5.735 1.85 5.905 2.36 ;
        RECT 4.495 1.68 5.905 1.85 ;
        RECT 4.495 1.45 4.825 1.68 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.14 1.015 1.31 ;
        RECT 0.125 1.31 0.355 1.48 ;
        RECT 0.685 1.11 1.015 1.14 ;
        RECT 0.125 1.48 0.895 1.65 ;
        RECT 0.685 0.94 2.015 1.11 ;
        RECT 0.565 1.65 0.895 1.78 ;
        RECT 0.685 0.35 1.015 0.94 ;
        RECT 1.685 0.35 2.015 0.94 ;
        RECT 0.565 1.78 1.895 1.95 ;
        RECT 0.565 1.95 0.895 2.98 ;
        RECT 1.565 1.95 1.895 2.98 ;
    END
    ANTENNADIFFAREA 1.3133 ;
  END X

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845 1.12 7.295 1.41 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.075 1.58 8.035 1.78 ;
        RECT 6.075 1.78 6.405 1.8 ;
        RECT 7.565 1.45 8.035 1.58 ;
        RECT 6.075 1.13 6.405 1.58 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.065 1.18 5.735 1.51 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A3

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.925 1.27 4.255 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.655 2.7 4.025 2.96 ;
      RECT 4.73 0.96 5.06 1.01 ;
      RECT 4.73 0.95 6.06 0.96 ;
      RECT 4.73 0.79 8.045 0.95 ;
      RECT 7.715 0.95 8.045 1.03 ;
      RECT 5.73 0.78 8.045 0.79 ;
      RECT 4.73 0.425 5.06 0.79 ;
      RECT 5.73 0.35 6.06 0.78 ;
      RECT 6.74 0.35 6.99 0.78 ;
      RECT 7.715 0.35 8.045 0.78 ;
      RECT 2.8 0.255 5.06 0.425 ;
      RECT 2.8 0.425 3.13 0.94 ;
      RECT 3.73 0.425 4.06 0.76 ;
      RECT 6.155 2.2 6.675 2.22 ;
      RECT 6.155 1.97 7.595 2.2 ;
      RECT 7.265 1.95 7.595 1.97 ;
      RECT 3.23 2.02 5.565 2.19 ;
      RECT 3.3 0.93 4.56 1.1 ;
      RECT 4.23 0.595 4.56 0.93 ;
      RECT 1.255 1.28 2.355 1.61 ;
      RECT 3.23 1.92 3.575 2.02 ;
      RECT 3.23 1.28 3.56 1.92 ;
      RECT 2.185 1.11 3.56 1.28 ;
      RECT 3.3 1.1 3.56 1.11 ;
      RECT 3.3 0.595 3.56 0.93 ;
      RECT 4.785 2.7 6.245 2.98 ;
      RECT 6.075 2.56 6.245 2.7 ;
      RECT 6.075 2.39 8.045 2.56 ;
      RECT 7.715 2.56 8.045 2.98 ;
      RECT 7.765 1.95 8.045 2.39 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 2.24 0.085 2.57 0.94 ;
      RECT 5.23 0.085 5.56 0.62 ;
      RECT 6.23 0.085 6.56 0.61 ;
      RECT 7.16 0.085 7.545 0.6 ;
      RECT 0.185 0.085 0.515 0.97 ;
      RECT 1.185 0.085 1.515 0.77 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 6.805 2.73 7.135 3.245 ;
      RECT 2.085 1.95 2.415 3.245 ;
      RECT 0.115 1.82 0.365 3.245 ;
      RECT 1.065 2.12 1.395 3.245 ;
      RECT 4.195 2.7 4.525 3.245 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
  END
END scs8ls_o32a_4

MACRO scs8ls_o32ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.88 1.18 3.235 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 2.445 2.89 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.35 1.875 2.52 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.18 0.445 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.975 1.35 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635 1.95 1.375 2.98 ;
        RECT 0.635 1.13 0.805 1.95 ;
        RECT 0.615 0.72 1.14 1.13 ;
    END
    ANTENNADIFFAREA 0.9929 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.115 0.35 1.68 0.52 ;
      RECT 1.35 0.52 1.68 1.01 ;
      RECT 1.35 1.01 2.71 1.18 ;
      RECT 2.38 0.35 2.71 1.01 ;
      RECT 0.115 0.52 0.445 1.01 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.835 1.82 3.165 3.245 ;
      RECT 0.135 1.82 0.465 3.245 ;
      RECT 1.85 0.085 2.18 0.81 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.88 0.085 3.14 1.01 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o32ai_1

MACRO scs8ls_o211a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.335 1.47 2.005 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325 0.255 3.715 0.64 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.49 3.335 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.635 1.49 4.195 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END C1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.82 0.445 2.98 ;
        RECT 0.085 1.13 0.255 1.82 ;
        RECT 0.085 0.35 0.445 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.265 1.13 2.495 1.3 ;
      RECT 2.325 0.98 2.495 1.13 ;
      RECT 1.265 0.66 1.595 1.13 ;
      RECT 2.325 0.81 3.185 0.98 ;
      RECT 0.925 1.97 4.205 2.14 ;
      RECT 3.875 2.14 4.205 2.98 ;
      RECT 2.665 1.15 4.135 1.32 ;
      RECT 3.76 0.835 4.135 1.15 ;
      RECT 3.885 0.66 4.135 0.835 ;
      RECT 2.395 2.14 2.725 2.98 ;
      RECT 2.395 1.94 2.835 1.97 ;
      RECT 2.665 1.32 2.835 1.94 ;
      RECT 0.925 1.65 1.095 1.97 ;
      RECT 0.425 1.32 1.095 1.65 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 0.615 0.085 0.945 1.13 ;
      RECT 1.765 0.085 2.155 0.925 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 0.615 2.31 1.855 3.245 ;
      RECT 2.895 2.31 3.705 3.245 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_o211a_1

MACRO scs8ls_o211a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.98 0.35 3.235 1.13 ;
        RECT 3.005 1.13 3.235 1.41 ;
        RECT 3.005 1.41 3.225 1.82 ;
        RECT 2.895 1.82 3.225 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.35 1.125 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965 1.35 2.295 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.435 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END C1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.335 1.35 1.795 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.025 0.67 2.35 0.84 ;
      RECT 1.025 0.35 1.355 0.67 ;
      RECT 2.02 0.35 2.35 0.67 ;
      RECT 0.105 1.95 2.675 2.12 ;
      RECT 2.505 1.63 2.675 1.95 ;
      RECT 2.505 1.3 2.835 1.63 ;
      RECT 2.505 1.18 2.675 1.3 ;
      RECT 0.605 1.01 2.675 1.18 ;
      RECT 1.105 2.12 1.435 2.86 ;
      RECT 0.13 0.35 0.775 1.01 ;
      RECT 0.105 2.12 0.435 2.86 ;
      RECT 0.105 1.82 0.435 1.95 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 3.395 1.82 3.725 3.245 ;
      RECT 0.605 2.29 0.935 3.245 ;
      RECT 2.025 2.29 2.725 3.245 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 3.41 0.085 3.74 1.13 ;
      RECT 1.525 0.085 1.775 0.5 ;
      RECT 2.55 0.085 2.8 0.84 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o211a_2

MACRO scs8ls_o211a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.13 0.355 1.8 ;
        RECT 0.125 1.8 1.945 1.97 ;
        RECT 0.125 0.96 1.76 1.13 ;
        RECT 0.615 1.97 0.945 2.98 ;
        RECT 1.615 1.97 1.945 2.98 ;
        RECT 0.58 0.35 0.83 0.96 ;
        RECT 1.51 0.35 1.76 0.96 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END X

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.45 1.45 3.78 1.78 ;
    END
    ANTENNAGATEAREA 0.444 ;
  END C1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505 1.435 2.835 1.78 ;
    END
    ANTENNAGATEAREA 0.444 ;
  END B1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.45 5.835 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.075 1.45 6.595 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.115 1.95 5.655 2.12 ;
      RECT 5.325 2.12 5.655 2.735 ;
      RECT 3.79 2.12 4.12 2.815 ;
      RECT 3.95 1.28 4.12 1.95 ;
      RECT 3.39 1.11 4.12 1.28 ;
      RECT 3.39 0.935 3.72 1.11 ;
      RECT 2.775 2.12 3.105 2.815 ;
      RECT 2.115 1.63 2.285 1.95 ;
      RECT 0.615 1.3 2.285 1.63 ;
      RECT 4.825 2.905 6.105 3.075 ;
      RECT 4.825 2.29 5.155 2.905 ;
      RECT 5.855 1.95 6.105 2.905 ;
      RECT 0 3.245 6.72 3.415 ;
      RECT 2.115 2.29 2.445 3.245 ;
      RECT 3.275 2.29 3.605 3.245 ;
      RECT 4.325 2.29 4.655 3.245 ;
      RECT 6.275 1.95 6.605 3.245 ;
      RECT 0.115 2.14 0.445 3.245 ;
      RECT 1.115 2.14 1.445 3.245 ;
      RECT 0 -0.085 6.72 0.085 ;
      RECT 1.94 0.085 2.27 1.13 ;
      RECT 4.83 0.085 5.175 0.935 ;
      RECT 5.775 0.085 6.105 0.94 ;
      RECT 0.15 0.085 0.4 0.79 ;
      RECT 1.01 0.085 1.34 0.79 ;
      RECT 3.04 0.765 3.21 1.285 ;
      RECT 3.04 0.595 4.22 0.765 ;
      RECT 3.89 0.765 4.22 0.94 ;
      RECT 4.4 1.28 4.65 1.285 ;
      RECT 4.4 1.11 6.605 1.28 ;
      RECT 5.345 0.605 5.595 1.11 ;
      RECT 6.275 0.605 6.605 1.11 ;
      RECT 4.4 0.425 4.65 1.11 ;
      RECT 2.53 0.255 4.65 0.425 ;
      RECT 2.53 0.425 2.78 1.265 ;
    LAYER mcon ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o211a_4

MACRO scs8ls_o211ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.3 0.435 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.63 0.835 2.89 ;
        RECT 0.605 1.55 1.165 1.63 ;
        RECT 0.665 1.3 1.165 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975 1.18 2.305 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END C1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 0.44 2.77 1.01 ;
        RECT 2.595 1.01 2.77 1.8 ;
        RECT 1.125 1.8 2.77 1.97 ;
        RECT 1.125 1.97 1.455 2.98 ;
        RECT 2.205 1.97 2.77 2.98 ;
    END
    ANTENNADIFFAREA 1.4276 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.44 1.795 1.3 ;
        RECT 1.405 1.3 1.795 1.63 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.135 0.96 1.395 1.13 ;
      RECT 0.135 0.35 0.465 0.96 ;
      RECT 1.145 0.35 1.395 0.96 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 0.115 1.95 0.365 3.245 ;
      RECT 1.705 2.14 2.035 3.245 ;
      RECT 0 -0.085 2.88 0.085 ;
      RECT 0.635 0.085 0.965 0.78 ;
    LAYER mcon ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o211ai_1

MACRO scs8ls_o211ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 2.12 0.925 2.98 ;
        RECT 0.595 1.95 3.285 2.12 ;
        RECT 1.495 2.12 1.825 2.98 ;
        RECT 2.955 2.12 3.285 2.735 ;
        RECT 0.72 1.18 0.89 1.95 ;
        RECT 0.56 0.595 0.89 1.18 ;
    END
    ANTENNADIFFAREA 1.2152 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.365 1.18 4.695 1.32 ;
        RECT 3.685 1.32 4.695 1.65 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.435 1.65 3.235 1.78 ;
        RECT 2.435 1.32 3.445 1.65 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.35 2.015 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 0.55 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END C1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.505 2.905 3.655 3.075 ;
      RECT 3.485 1.99 3.655 2.905 ;
      RECT 3.485 1.82 4.685 1.99 ;
      RECT 4.355 1.99 4.685 2.98 ;
      RECT 2.505 2.29 2.755 2.905 ;
      RECT 1.56 1.15 1.89 1.18 ;
      RECT 1.56 0.98 4.16 1.15 ;
      RECT 1.56 0.9 1.89 0.98 ;
      RECT 3.07 0.35 3.24 0.98 ;
      RECT 3.935 0.35 4.16 0.98 ;
      RECT 1.06 0.73 1.39 1.18 ;
      RECT 1.06 0.425 2.33 0.73 ;
      RECT 0.13 0.255 2.33 0.425 ;
      RECT 0.13 0.425 0.38 1.18 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 3.855 2.16 4.185 3.245 ;
      RECT 0.145 1.95 0.395 3.245 ;
      RECT 1.125 2.29 1.295 3.245 ;
      RECT 2.025 2.29 2.275 3.245 ;
      RECT 2.56 0.085 2.89 0.795 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 3.42 0.085 3.75 0.795 ;
      RECT 4.33 0.085 4.685 1.01 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o211ai_2

MACRO scs8ls_o211ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.365 1.55 8.035 1.95 ;
        RECT 2.43 1.95 8.035 2.12 ;
        RECT 7.365 1.18 7.545 1.55 ;
        RECT 7.545 2.12 8.035 2.89 ;
        RECT 2.43 2.12 2.76 2.735 ;
        RECT 3.38 2.12 3.71 2.735 ;
        RECT 4.94 2.12 5.27 2.98 ;
        RECT 5.94 2.12 6.27 2.98 ;
        RECT 6.505 1.01 7.545 1.18 ;
        RECT 6.505 0.595 6.675 1.01 ;
        RECT 7.365 0.595 7.545 1.01 ;
    END
    ANTENNADIFFAREA 1.9152 ;
  END Y

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.87 1.35 7.075 1.78 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END C1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.35 5.635 1.78 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END B1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 4.195 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.795 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.115 1.01 5.765 1.18 ;
      RECT 3.795 0.82 4.905 1.01 ;
      RECT 5.435 0.595 5.765 1.01 ;
      RECT 0.115 0.35 0.445 1.01 ;
      RECT 1.125 0.35 1.375 1.01 ;
      RECT 2.055 0.35 2.225 1.01 ;
      RECT 2.915 0.35 3.085 1.01 ;
      RECT 3.795 0.35 3.965 0.82 ;
      RECT 4.145 0.255 8.045 0.425 ;
      RECT 7.715 0.425 8.045 1.18 ;
      RECT 5.085 0.65 5.255 0.84 ;
      RECT 4.145 0.425 5.255 0.65 ;
      RECT 5.995 0.425 6.325 1.18 ;
      RECT 6.855 0.425 7.185 0.84 ;
      RECT 1.93 2.905 4.21 3.075 ;
      RECT 3.88 2.29 4.21 2.905 ;
      RECT 1.93 2.12 2.26 2.905 ;
      RECT 0.13 1.95 2.26 2.12 ;
      RECT 0.13 2.12 0.46 2.98 ;
      RECT 1.03 2.12 1.36 2.98 ;
      RECT 2.96 2.29 3.21 2.905 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 0.66 2.29 0.83 3.245 ;
      RECT 1.56 2.29 1.73 3.245 ;
      RECT 4.44 2.29 4.77 3.245 ;
      RECT 5.44 2.29 5.77 3.245 ;
      RECT 6.44 2.29 7.29 3.245 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 0.615 0.085 0.945 0.84 ;
      RECT 1.545 0.085 1.875 0.84 ;
      RECT 2.405 0.085 2.735 0.84 ;
      RECT 3.265 0.085 3.595 0.84 ;
    LAYER mcon ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
  END
END scs8ls_o211ai_4

MACRO scs8ls_o21a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.3 2.775 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.445 1.435 1.78 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END B1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.715 1.445 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.35 0.365 1.82 ;
        RECT 0.115 1.82 0.445 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.575 0.96 2.765 1.13 ;
      RECT 1.575 0.35 1.825 0.96 ;
      RECT 2.515 0.35 2.765 0.96 ;
      RECT 1.36 2.12 1.69 2.795 ;
      RECT 0.695 1.95 1.69 2.12 ;
      RECT 0.535 1.105 1.395 1.275 ;
      RECT 1.145 0.35 1.395 1.105 ;
      RECT 0.695 1.55 0.865 1.95 ;
      RECT 0.535 1.275 0.865 1.55 ;
      RECT 0.545 0.085 0.875 0.935 ;
      RECT 0 -0.085 2.88 0.085 ;
      RECT 2.005 0.085 2.335 0.79 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 0.615 2.29 1.18 3.245 ;
      RECT 2.435 1.95 2.765 3.245 ;
    LAYER mcon ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_o21a_1

MACRO scs8ls_o21a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.965 0.35 3.295 1.72 ;
        RECT 2.465 1.72 3.295 1.89 ;
        RECT 2.465 1.89 2.795 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.18 1.955 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055 1.18 1.385 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.835 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.25 0.84 1.735 1.01 ;
      RECT 0.25 0.34 0.58 0.84 ;
      RECT 1.405 0.34 1.735 0.84 ;
      RECT 2.125 1.22 2.645 1.55 ;
      RECT 1.325 1.89 1.655 2.86 ;
      RECT 1.325 1.72 2.295 1.89 ;
      RECT 2.125 1.55 2.295 1.72 ;
      RECT 2.125 1.01 2.295 1.22 ;
      RECT 1.905 0.34 2.295 1.01 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 2.965 2.06 3.295 3.245 ;
      RECT 1.965 2.06 2.295 3.245 ;
      RECT 0.335 1.82 0.665 3.245 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 3.475 0.085 3.725 1.13 ;
      RECT 0.75 0.085 1.235 0.6 ;
      RECT 2.465 0.085 2.795 1.05 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o21a_2

MACRO scs8ls_o21a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.965 1.55 5.635 1.72 ;
        RECT 3.815 1.72 5.635 1.78 ;
        RECT 4.965 1.005 5.135 1.55 ;
        RECT 3.815 1.78 5.145 1.89 ;
        RECT 3.99 0.835 5.135 1.005 ;
        RECT 3.815 1.89 4.145 2.98 ;
        RECT 4.815 1.89 5.145 2.98 ;
        RECT 4.965 0.35 5.135 0.835 ;
        RECT 3.99 0.33 4.24 0.835 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END X

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.515 3.235 1.78 ;
    END
    ANTENNAGATEAREA 0.444 ;
  END B1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835 1.445 1.505 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.795 1.445 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.615 2.905 1.895 3.075 ;
      RECT 1.565 2.29 1.895 2.905 ;
      RECT 0.615 1.95 0.865 2.905 ;
      RECT 0.115 1.275 0.445 1.285 ;
      RECT 0.115 1.105 2.39 1.275 ;
      RECT 0.115 0.605 0.445 1.105 ;
      RECT 1.13 0.605 1.38 1.105 ;
      RECT 2.06 0.435 2.39 1.105 ;
      RECT 2.06 0.265 3.33 0.435 ;
      RECT 3 0.435 3.33 1.005 ;
      RECT 3.405 1.345 4.795 1.55 ;
      RECT 2.57 1.175 4.795 1.345 ;
      RECT 1.065 1.95 3.575 2.12 ;
      RECT 2.565 2.12 2.895 2.795 ;
      RECT 3.405 1.55 3.575 1.95 ;
      RECT 2.57 0.605 2.82 1.175 ;
      RECT 1.065 2.12 1.395 2.735 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 5.315 1.95 5.645 3.245 ;
      RECT 3.135 2.3 3.615 3.245 ;
      RECT 2.065 2.29 2.395 3.245 ;
      RECT 0.115 1.915 0.445 3.245 ;
      RECT 4.315 2.06 4.645 3.245 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 5.315 0.085 5.645 1.13 ;
      RECT 0.615 0.085 0.95 0.935 ;
      RECT 1.56 0.085 1.89 0.935 ;
      RECT 3.56 0.085 3.81 1.005 ;
      RECT 4.42 0.085 4.785 0.665 ;
    LAYER mcon ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o21a_4

MACRO scs8ls_o21ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.555 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.35 1.395 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.35 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.725 1.95 1.545 2.98 ;
        RECT 0.725 1.18 0.895 1.95 ;
        RECT 0.725 1.01 2.285 1.18 ;
        RECT 1.955 0.35 2.285 1.01 ;
    END
    ANTENNADIFFAREA 0.8283 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.115 0.84 0.445 1.01 ;
      RECT 0.115 0.67 1.785 0.84 ;
      RECT 0.115 0.35 0.42 0.67 ;
      RECT 1.48 0.35 1.785 0.67 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 0.605 0.085 1.295 0.5 ;
      RECT 0 3.245 2.4 3.415 ;
      RECT 1.87 1.95 2.2 3.245 ;
      RECT 0.305 1.82 0.555 3.245 ;
    LAYER mcon ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_o21ai_1

MACRO scs8ls_o21ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.82 2.795 2.29 ;
        RECT 1.065 2.29 2.795 2.46 ;
        RECT 2.525 1.13 2.735 1.82 ;
        RECT 2.525 2.46 2.795 2.98 ;
        RECT 1.065 2.46 1.395 2.735 ;
        RECT 2.475 0.715 2.735 1.13 ;
    END
    ANTENNADIFFAREA 0.9611 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.755 1.35 2.275 1.95 ;
        RECT 0.265 1.95 2.275 2.12 ;
        RECT 0.265 1.35 0.595 1.95 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.845 1.35 1.515 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.18 3.235 1.55 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.565 2.905 1.895 3.075 ;
      RECT 1.565 2.63 1.895 2.905 ;
      RECT 0.565 2.29 0.895 2.905 ;
      RECT 2.055 0.35 3.245 0.52 ;
      RECT 2.915 0.52 3.245 1.01 ;
      RECT 0.115 1.01 2.305 1.18 ;
      RECT 2.055 0.52 2.305 1.01 ;
      RECT 0.115 0.35 0.445 1.01 ;
      RECT 1.125 0.35 1.375 1.01 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.995 1.82 3.245 3.245 ;
      RECT 2.095 2.63 2.345 3.245 ;
      RECT 0.115 2.29 0.365 3.245 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 0.615 0.085 0.945 0.83 ;
      RECT 1.545 0.085 1.875 0.83 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o21ai_2

MACRO scs8ls_o21ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.18 3.165 1.55 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END B1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.35 5.635 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.65 1.795 1.78 ;
        RECT 0.445 1.32 1.795 1.65 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.335 1.55 3.715 1.82 ;
        RECT 2.365 1.82 3.715 1.95 ;
        RECT 3.335 1.01 3.505 1.55 ;
        RECT 2.365 1.95 5.19 2.12 ;
        RECT 2.28 0.84 3.505 1.01 ;
        RECT 3.96 2.12 4.29 2.735 ;
        RECT 4.86 2.12 5.19 2.735 ;
        RECT 2.28 0.595 2.53 0.84 ;
        RECT 3.22 0.595 3.505 0.84 ;
    END
    ANTENNADIFFAREA 1.4784 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 4.025 0.085 4.355 0.84 ;
      RECT 4.885 0.085 5.215 0.84 ;
      RECT 0.545 0.085 0.875 0.81 ;
      RECT 1.405 0.085 1.735 0.67 ;
      RECT 1.93 0.255 3.845 0.425 ;
      RECT 3.675 0.425 3.845 1.01 ;
      RECT 3.675 1.01 5.645 1.18 ;
      RECT 4.535 0.35 4.705 1.01 ;
      RECT 5.395 0.35 5.645 1.01 ;
      RECT 0.115 1.01 1.225 1.15 ;
      RECT 0.115 0.98 2.1 1.01 ;
      RECT 1.055 0.84 2.1 0.98 ;
      RECT 0.115 0.35 0.365 0.98 ;
      RECT 1.93 0.425 2.1 0.84 ;
      RECT 1.055 0.35 1.225 0.84 ;
      RECT 2.71 0.425 3.04 0.67 ;
      RECT 3.46 2.905 5.64 3.075 ;
      RECT 5.39 1.95 5.64 2.905 ;
      RECT 1.465 2.46 1.795 2.98 ;
      RECT 1.465 2.12 1.795 2.29 ;
      RECT 0.565 1.95 1.795 2.12 ;
      RECT 0.565 2.12 0.895 2.98 ;
      RECT 0.565 1.82 0.895 1.95 ;
      RECT 1.465 2.29 3.79 2.46 ;
      RECT 3.46 2.46 3.79 2.905 ;
      RECT 4.49 2.29 4.66 2.905 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 1.995 2.63 2.245 3.245 ;
      RECT 1.095 2.29 1.265 3.245 ;
      RECT 0.115 1.82 0.365 3.245 ;
      RECT 2.9 2.63 3.23 3.245 ;
    LAYER mcon ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o21ai_4

MACRO scs8ls_o21ba_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395 1.82 3.755 2.98 ;
        RECT 3.585 1.13 3.755 1.82 ;
        RECT 3.39 0.35 3.755 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.13 0.55 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835 1.13 1.315 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.515 1.18 2.845 1.55 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END B1N

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.115 0.79 1.445 0.96 ;
      RECT 0.115 0.35 0.445 0.79 ;
      RECT 1.115 0.35 1.445 0.79 ;
      RECT 1.975 1.82 2.69 2.15 ;
      RECT 2.135 0.68 2.72 1.01 ;
      RECT 1.975 1.22 2.305 1.82 ;
      RECT 2.135 1.01 2.305 1.22 ;
      RECT 3.055 1.32 3.415 1.65 ;
      RECT 1.055 2.32 3.225 2.49 ;
      RECT 3.055 1.65 3.225 2.32 ;
      RECT 1.055 2.49 1.385 2.98 ;
      RECT 1.055 1.97 1.785 2.32 ;
      RECT 1.615 1.03 1.785 1.97 ;
      RECT 1.615 0.35 1.945 1.03 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 0.615 0.085 0.945 0.62 ;
      RECT 2.89 0.085 3.22 1.01 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 1.555 2.66 1.885 3.245 ;
      RECT 2.895 2.66 3.225 3.245 ;
      RECT 0.115 1.97 0.445 3.245 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_o21ba_1

MACRO scs8ls_o21ba_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.3 0.455 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END B1N

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.72 1.18 3.235 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.01 0.35 1.34 1.13 ;
        RECT 1.01 1.13 1.18 1.82 ;
        RECT 1.01 1.82 1.44 2.07 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.18 3.735 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.41 0.84 3.74 1.01 ;
      RECT 2.41 0.67 3.74 0.84 ;
      RECT 2.41 0.35 2.74 0.67 ;
      RECT 3.41 0.35 3.74 0.67 ;
      RECT 2.445 2.41 2.775 2.86 ;
      RECT 2.38 1.82 2.775 2.41 ;
      RECT 2.38 1.18 2.55 1.82 ;
      RECT 1.51 1.01 2.55 1.18 ;
      RECT 1.51 1.18 1.68 1.3 ;
      RECT 1.98 0.35 2.23 1.01 ;
      RECT 1.35 1.3 1.68 1.63 ;
      RECT 0.115 2.24 2.21 2.41 ;
      RECT 1.89 1.35 2.21 2.24 ;
      RECT 0.115 2.41 0.445 2.7 ;
      RECT 0.115 1.95 0.795 2.24 ;
      RECT 0.625 1.13 0.795 1.95 ;
      RECT 0.105 0.96 0.795 1.13 ;
      RECT 0.105 0.455 0.355 0.96 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 1.565 2.58 2.235 3.245 ;
      RECT 3.405 1.82 3.735 3.245 ;
      RECT 0.65 2.58 0.98 3.245 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 1.52 0.085 1.77 0.82 ;
      RECT 2.91 0.085 3.24 0.5 ;
      RECT 0.535 0.085 0.785 0.79 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o21ba_2

MACRO scs8ls_o21ba_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.55 1.315 1.82 ;
        RECT 1.085 1.82 2.345 2.22 ;
        RECT 1.145 1.12 1.315 1.55 ;
        RECT 1.145 0.95 2.21 1.12 ;
        RECT 1.145 0.35 1.34 0.95 ;
        RECT 1.96 0.35 2.21 0.95 ;
    END
    ANTENNADIFFAREA 1.0938 ;
  END X

  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.18 0.835 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1N

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.845 1.45 6.115 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175 1.45 4.675 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.085 2.39 3.32 2.56 ;
      RECT 3.15 1.96 3.32 2.39 ;
      RECT 3.15 1.63 3.49 1.96 ;
      RECT 0.085 2.56 0.445 2.98 ;
      RECT 0.085 1.82 0.445 2.39 ;
      RECT 0.085 0.35 0.475 1.01 ;
      RECT 0.085 1.01 0.255 1.82 ;
      RECT 0 3.245 6.24 3.415 ;
      RECT 1.565 2.73 1.895 3.245 ;
      RECT 2.465 2.73 3.205 3.245 ;
      RECT 3.945 2.47 4.275 3.245 ;
      RECT 5.875 1.95 6.125 3.245 ;
      RECT 0.615 2.73 0.995 3.245 ;
      RECT 0 -0.085 6.24 0.085 ;
      RECT 2.39 0.085 2.64 1.12 ;
      RECT 4.5 0.085 4.75 0.94 ;
      RECT 5.36 0.085 5.61 0.94 ;
      RECT 0.645 0.085 0.975 1.01 ;
      RECT 1.53 0.085 1.78 0.78 ;
      RECT 4.445 2.905 5.675 3.075 ;
      RECT 4.445 2.47 4.775 2.905 ;
      RECT 5.345 1.95 5.675 2.905 ;
      RECT 4 1.12 6.125 1.28 ;
      RECT 3.15 1.11 6.125 1.12 ;
      RECT 3.15 0.95 4.33 1.11 ;
      RECT 4.93 0.605 5.18 1.11 ;
      RECT 5.79 0.605 6.125 1.11 ;
      RECT 4 0.605 4.33 0.95 ;
      RECT 3.15 0.595 3.32 0.95 ;
      RECT 3.49 2.13 5.145 2.3 ;
      RECT 4.975 2.3 5.145 2.735 ;
      RECT 3.66 1.95 5.145 2.13 ;
      RECT 3.49 2.3 3.74 2.98 ;
      RECT 3.66 1.46 3.83 1.95 ;
      RECT 1.485 1.29 3.83 1.46 ;
      RECT 1.485 1.46 2.98 1.62 ;
      RECT 2.81 0.425 2.98 1.29 ;
      RECT 2.81 0.255 3.83 0.425 ;
      RECT 3.5 0.425 3.83 0.78 ;
    LAYER mcon ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o21ba_4

MACRO scs8ls_o21bai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.3 2.775 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.63 2.275 2.89 ;
        RECT 1.75 1.3 2.275 1.63 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475 1.99 1.84 2.98 ;
        RECT 1.305 1.82 1.84 1.99 ;
        RECT 1.305 1.13 1.475 1.82 ;
        RECT 1.085 0.35 1.475 1.13 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END Y

  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.45 0.565 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END B1N

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.645 0.96 2.765 1.13 ;
      RECT 1.645 0.35 1.815 0.96 ;
      RECT 2.515 0.35 2.765 0.96 ;
      RECT 0.745 1.3 1.135 1.63 ;
      RECT 0.135 2.12 0.465 2.98 ;
      RECT 0.135 1.95 0.915 2.12 ;
      RECT 0.745 1.63 0.915 1.95 ;
      RECT 0.745 1.28 0.915 1.3 ;
      RECT 0.11 1.11 0.915 1.28 ;
      RECT 0.11 0.35 0.36 1.11 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 2.52 1.95 2.77 3.245 ;
      RECT 0.635 2.29 1.305 3.245 ;
      RECT 0 -0.085 2.88 0.085 ;
      RECT 1.995 0.085 2.335 0.68 ;
      RECT 0.54 0.085 0.87 0.94 ;
    LAYER mcon ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o21bai_1

MACRO scs8ls_o21bai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.53 1.18 1.865 2.29 ;
        RECT 1.53 2.29 3.22 2.46 ;
        RECT 1.615 0.615 1.865 1.18 ;
        RECT 1.53 2.46 1.78 2.98 ;
        RECT 3.05 2.46 3.22 2.735 ;
    END
    ANTENNADIFFAREA 0.8792 ;
  END Y

  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.46 1.35 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1N

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.82 1.35 3.235 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.65 3.715 1.95 ;
        RECT 3.485 1.32 4.055 1.65 ;
        RECT 2.25 1.95 3.715 2.12 ;
        RECT 2.25 1.35 2.58 1.95 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.035 1.15 3.245 1.18 ;
      RECT 2.035 1.01 4.185 1.15 ;
      RECT 3.075 0.98 4.185 1.01 ;
      RECT 2.035 0.425 2.365 1.01 ;
      RECT 3.075 0.35 3.245 0.98 ;
      RECT 3.935 0.35 4.185 0.98 ;
      RECT 1.105 0.255 2.365 0.425 ;
      RECT 1.105 0.425 1.435 0.84 ;
      RECT 2.52 2.905 3.755 3.075 ;
      RECT 3.42 2.29 3.755 2.905 ;
      RECT 2.52 2.63 2.85 2.905 ;
      RECT 0.115 1.95 0.64 2.86 ;
      RECT 0.115 1.01 1.36 1.18 ;
      RECT 1.03 1.18 1.36 1.55 ;
      RECT 0.115 1.18 0.285 1.95 ;
      RECT 0.115 0.35 0.365 1.01 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 3.955 1.82 4.205 3.245 ;
      RECT 1.005 1.82 1.335 3.245 ;
      RECT 1.98 2.65 2.35 3.245 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 2.535 0.085 2.865 0.84 ;
      RECT 3.425 0.085 3.755 0.81 ;
      RECT 0.545 0.085 0.875 0.84 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o21bai_2

MACRO scs8ls_o21bai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.45 7.075 1.78 ;
    END
    ANTENNAGATEAREA 0.363 ;
  END B1N

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.35 3.715 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.795 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.18 4.195 1.95 ;
        RECT 2.37 1.95 5.625 2.02 ;
        RECT 3.965 1.01 5.595 1.18 ;
        RECT 2.37 2.02 4.71 2.12 ;
        RECT 5.295 2.02 5.625 2.98 ;
        RECT 4.38 1.85 5.625 1.95 ;
        RECT 4.265 0.595 4.595 1.01 ;
        RECT 5.265 0.595 5.595 1.01 ;
        RECT 2.37 2.12 2.62 2.735 ;
        RECT 3.32 2.12 3.65 2.735 ;
        RECT 4.38 2.12 4.71 2.98 ;
    END
    ANTENNADIFFAREA 1.855 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.765 0.255 6.095 0.425 ;
      RECT 5.765 0.425 6.095 0.94 ;
      RECT 0.115 1.01 3.075 1.18 ;
      RECT 2.825 0.84 3.075 1.01 ;
      RECT 0.115 0.35 0.365 1.01 ;
      RECT 1.105 0.35 1.275 1.01 ;
      RECT 1.965 0.35 2.135 1.01 ;
      RECT 2.825 0.35 3.075 0.67 ;
      RECT 2.825 0.67 4.095 0.84 ;
      RECT 3.765 0.425 4.095 0.67 ;
      RECT 4.765 0.425 5.095 0.84 ;
      RECT 6.305 2.12 6.555 2.98 ;
      RECT 5.795 1.95 6.555 2.12 ;
      RECT 5.795 1.11 6.575 1.28 ;
      RECT 6.325 0.5 6.575 1.11 ;
      RECT 5.795 1.68 5.965 1.95 ;
      RECT 4.37 1.35 5.965 1.68 ;
      RECT 5.795 1.28 5.965 1.35 ;
      RECT 2 2.905 4.15 3.075 ;
      RECT 3.82 2.29 4.15 2.905 ;
      RECT 2 2.12 2.17 2.905 ;
      RECT 0.12 1.95 2.17 2.12 ;
      RECT 0.12 2.12 0.37 2.98 ;
      RECT 1.02 2.12 1.27 2.98 ;
      RECT 2 1.82 2.17 1.95 ;
      RECT 2.82 2.29 3.15 2.905 ;
      RECT 0 3.245 7.2 3.415 ;
      RECT 5.855 2.29 6.105 3.245 ;
      RECT 6.755 2.1 7.085 3.245 ;
      RECT 0.57 2.29 0.82 3.245 ;
      RECT 1.47 2.29 1.8 3.245 ;
      RECT 4.91 2.19 5.08 3.245 ;
      RECT 0 -0.085 7.2 0.085 ;
      RECT 6.755 0.085 7.085 1.28 ;
      RECT 0.545 0.085 0.875 0.84 ;
      RECT 1.455 0.085 1.785 0.84 ;
      RECT 2.315 0.085 2.645 0.84 ;
      RECT 3.255 0.085 3.585 0.5 ;
    LAYER mcon ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
  END
END scs8ls_o21bai_4

MACRO scs8ls_o221a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.35 0.52 1.13 ;
        RECT 0.115 1.13 0.285 1.82 ;
        RECT 0.115 1.82 0.445 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.145 1.45 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.46 3.255 1.79 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.45 1.905 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.45 1.335 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.12 3.825 1.79 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END C1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.26 0.425 2.59 0.94 ;
      RECT 2.26 0.255 3.6 0.425 ;
      RECT 3.27 0.425 3.6 0.95 ;
      RECT 1.2 1.11 3.1 1.28 ;
      RECT 2.77 0.595 3.1 1.11 ;
      RECT 1.2 0.45 1.53 1.11 ;
      RECT 1.725 2.12 4.205 2.13 ;
      RECT 3.875 2.13 4.205 2.98 ;
      RECT 0.615 1.96 4.205 2.12 ;
      RECT 4.035 0.95 4.205 1.96 ;
      RECT 3.77 0.36 4.205 0.95 ;
      RECT 1.725 2.13 2.055 2.98 ;
      RECT 0.615 1.95 2.055 1.96 ;
      RECT 0.615 1.65 0.785 1.95 ;
      RECT 0.455 1.32 0.785 1.65 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 2.865 2.3 3.705 3.245 ;
      RECT 0.68 2.29 1.06 3.245 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 0.69 0.085 1.02 1.13 ;
      RECT 1.7 0.085 2.03 0.94 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o221a_1

MACRO scs8ls_o221a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.35 1.395 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.79 0.35 4.265 1.13 ;
        RECT 4.095 1.13 4.265 1.82 ;
        RECT 3.905 1.82 4.265 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.435 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END C1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.35 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B2

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.485 1.35 2.815 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.35 3.385 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.945 0.52 1.115 1.13 ;
      RECT 0.945 0.35 2.13 0.52 ;
      RECT 1.8 0.52 2.13 0.83 ;
      RECT 1.295 1.01 3.12 1.18 ;
      RECT 1.295 0.8 1.62 1.01 ;
      RECT 2.87 0.35 3.12 1.01 ;
      RECT 3.565 1.32 3.925 1.65 ;
      RECT 0.115 1.95 3.735 2.12 ;
      RECT 3.565 1.65 3.735 1.95 ;
      RECT 2.065 2.12 2.395 2.86 ;
      RECT 0.115 2.12 0.445 2.86 ;
      RECT 0.115 1.82 0.775 1.95 ;
      RECT 0.605 1.01 0.775 1.82 ;
      RECT 0.37 0.35 0.775 1.01 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 4.435 1.82 4.685 3.245 ;
      RECT 0.615 2.29 1.525 3.245 ;
      RECT 3.405 2.29 3.735 3.245 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 4.435 0.085 4.685 1.13 ;
      RECT 2.36 0.085 2.69 0.83 ;
      RECT 3.29 0.085 3.62 1.13 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o221a_2

MACRO scs8ls_o221a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.445 0.89 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END C1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.445 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.445 4.195 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.365 1.445 4.695 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.35 5.32 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.785 1.55 7.555 1.78 ;
        RECT 6.785 1.78 7.115 1.85 ;
        RECT 6.785 1.18 7.065 1.55 ;
        RECT 5.83 1.85 7.115 2.02 ;
        RECT 5.735 1.01 7.065 1.18 ;
        RECT 5.83 2.02 6.16 2.98 ;
        RECT 6.785 2.02 7.115 2.98 ;
        RECT 5.735 0.475 5.985 1.01 ;
        RECT 6.735 0.475 7.065 1.01 ;
    END
    ANTENNADIFFAREA 1.2357 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.475 1.275 1.805 1.285 ;
      RECT 1.475 1.18 4.115 1.275 ;
      RECT 1.475 1.105 5.055 1.18 ;
      RECT 1.475 1.025 2.74 1.105 ;
      RECT 3.94 1.01 5.055 1.105 ;
      RECT 2.475 0.635 2.67 1.025 ;
      RECT 1.475 0.605 1.805 1.025 ;
      RECT 4.805 0.59 5.055 1.01 ;
      RECT 3.94 0.585 4.115 1.01 ;
      RECT 1.975 0.455 2.305 0.855 ;
      RECT 1.975 0.435 3.17 0.455 ;
      RECT 2.84 0.455 3.17 0.855 ;
      RECT 0.115 0.285 3.17 0.435 ;
      RECT 0.115 0.435 0.365 1.275 ;
      RECT 0.975 0.435 1.305 0.935 ;
      RECT 0.115 0.265 2.305 0.285 ;
      RECT 1.515 2.905 2.745 3.075 ;
      RECT 1.515 2.29 1.845 2.905 ;
      RECT 2.415 2.29 2.745 2.905 ;
      RECT 3.8 2.905 5.13 3.075 ;
      RECT 3.8 2.29 4.13 2.905 ;
      RECT 4.8 2.29 5.13 2.905 ;
      RECT 5.49 1.35 6.615 1.68 ;
      RECT 0.565 1.95 5.66 2.12 ;
      RECT 5.49 1.68 5.66 1.95 ;
      RECT 4.3 2.12 4.63 2.735 ;
      RECT 2.045 2.12 2.215 2.735 ;
      RECT 0.565 2.12 0.895 2.955 ;
      RECT 1.06 1.275 1.23 1.95 ;
      RECT 0.545 1.105 1.23 1.275 ;
      RECT 0.545 0.605 0.795 1.105 ;
      RECT 0 3.245 7.68 3.415 ;
      RECT 7.315 1.95 7.565 3.245 ;
      RECT 1.095 2.29 1.345 3.245 ;
      RECT 2.915 2.29 3.63 3.245 ;
      RECT 5.3 2.29 5.63 3.245 ;
      RECT 0.115 1.95 0.365 3.245 ;
      RECT 6.36 2.19 6.61 3.245 ;
      RECT 0 -0.085 7.68 0.085 ;
      RECT 7.235 0.085 7.565 1.255 ;
      RECT 3.43 0.085 3.76 0.935 ;
      RECT 4.295 0.085 4.625 0.84 ;
      RECT 5.235 0.085 5.565 1.18 ;
      RECT 6.165 0.085 6.565 0.805 ;
    LAYER mcon ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
  END
END scs8ls_o221a_4

MACRO scs8ls_o221ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.35 2.775 1.68 ;
        RECT 2.525 1.68 2.775 2.89 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.875 1.35 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.3 0.435 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END C1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.3 3.715 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.35 1.635 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.35 0.445 0.96 ;
        RECT 0.115 0.96 0.775 1.13 ;
        RECT 0.605 1.13 0.775 1.95 ;
        RECT 0.325 1.95 2.355 2.12 ;
        RECT 0.325 2.12 0.575 2.98 ;
        RECT 2.025 2.12 2.355 2.98 ;
    END
    ANTENNADIFFAREA 1.0117 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.615 0.52 0.945 0.77 ;
      RECT 0.615 0.35 2.005 0.52 ;
      RECT 1.675 0.52 2.005 0.795 ;
      RECT 1.175 1.13 2.505 1.18 ;
      RECT 1.175 1.01 3.725 1.13 ;
      RECT 1.175 0.8 1.505 1.01 ;
      RECT 2.175 0.96 3.725 1.01 ;
      RECT 2.175 0.35 2.505 0.96 ;
      RECT 3.395 0.35 3.725 0.96 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 3.165 1.95 3.495 3.245 ;
      RECT 0.745 2.29 1.56 3.245 ;
      RECT 2.675 0.085 3.225 0.79 ;
      RECT 0 -0.085 3.84 0.085 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o221ai_1

MACRO scs8ls_o221ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.345 1.35 4.675 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.52 1.35 2.85 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.3 0.435 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END C1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.35 5.635 1.95 ;
        RECT 3.645 1.95 5.635 2.12 ;
        RECT 3.645 1.35 3.975 1.95 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.35 2.275 1.95 ;
        RECT 1.085 1.95 3.405 2.12 ;
        RECT 3.075 1.35 3.405 1.95 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.595 0.875 2.29 ;
        RECT 0.605 2.29 4.615 2.46 ;
        RECT 0.605 2.46 0.855 2.98 ;
        RECT 2.365 2.46 2.695 2.735 ;
        RECT 4.365 2.46 4.615 2.735 ;
    END
    ANTENNADIFFAREA 1.232 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.055 1.01 3.28 1.18 ;
      RECT 2.045 0.595 2.215 1.01 ;
      RECT 2.895 0.595 3.28 1.01 ;
      RECT 1.055 0.425 1.305 1.01 ;
      RECT 0.115 0.255 1.305 0.425 ;
      RECT 0.115 0.425 0.365 1.13 ;
      RECT 1.865 2.905 3.195 3.075 ;
      RECT 2.865 2.63 3.195 2.905 ;
      RECT 1.865 2.63 2.195 2.905 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 5.315 2.29 5.645 3.245 ;
      RECT 0.155 1.95 0.405 3.245 ;
      RECT 1.055 2.63 1.695 3.245 ;
      RECT 3.365 2.63 3.695 3.245 ;
      RECT 3.88 0.085 4.21 0.82 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 4.88 0.085 5.21 0.82 ;
      RECT 3.865 2.905 5.145 3.075 ;
      RECT 4.815 2.29 5.145 2.905 ;
      RECT 3.865 2.63 4.195 2.905 ;
      RECT 3.46 1.01 5.645 1.18 ;
      RECT 3.46 0.425 3.71 1.01 ;
      RECT 4.38 0.405 4.71 1.01 ;
      RECT 5.39 0.405 5.645 1.01 ;
      RECT 1.535 0.255 3.71 0.425 ;
      RECT 1.535 0.425 1.865 0.82 ;
      RECT 2.395 0.425 2.725 0.82 ;
    LAYER mcon ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o221ai_2

MACRO scs8ls_o221ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285 1.26 9.955 1.78 ;
        RECT 6.405 1.09 8.455 1.26 ;
        RECT 6.21 1.26 6.575 1.59 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845 2.22 7.26 2.52 ;
        RECT 6.93 2.52 7.26 2.735 ;
        RECT 1.575 2.12 7.26 2.22 ;
        RECT 1.575 2.22 1.825 2.98 ;
        RECT 4.055 2.22 4.225 2.735 ;
        RECT 4.925 2.22 5.255 2.735 ;
        RECT 0.565 2.05 8.16 2.12 ;
        RECT 0.565 2.12 0.895 2.98 ;
        RECT 7.83 2.12 8.16 2.735 ;
        RECT 0.565 1.95 1.825 2.05 ;
        RECT 6.845 1.95 8.16 2.05 ;
        RECT 1.575 1.82 1.825 1.95 ;
        RECT 1.575 1.18 1.745 1.82 ;
        RECT 0.545 1.01 1.745 1.18 ;
        RECT 0.545 0.595 0.875 1.01 ;
        RECT 1.405 0.595 1.745 1.01 ;
    END
    ANTENNADIFFAREA 2.5144 ;
  END Y

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.185 1.18 5.195 1.54 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.405 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END C1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845 1.43 8.035 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405 1.35 6 1.71 ;
        RECT 2.545 1.71 6 1.88 ;
        RECT 2.545 1.35 3.555 1.71 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.915 1.01 4.015 1.18 ;
      RECT 1.915 0.77 3.155 1.01 ;
      RECT 3.685 0.77 5.735 1.01 ;
      RECT 1.915 0.425 2.165 0.77 ;
      RECT 5.405 1.01 5.735 1.05 ;
      RECT 0.115 0.255 2.165 0.425 ;
      RECT 0.115 0.425 0.375 1.18 ;
      RECT 1.045 0.425 1.235 0.84 ;
      RECT 3.525 2.905 5.755 3.075 ;
      RECT 5.425 2.39 5.755 2.905 ;
      RECT 2.525 2.56 2.855 2.98 ;
      RECT 2.525 2.39 3.855 2.56 ;
      RECT 3.525 2.56 3.855 2.905 ;
      RECT 4.425 2.39 4.755 2.905 ;
      RECT 6.425 2.905 8.53 3.075 ;
      RECT 8.36 2.12 8.53 2.905 ;
      RECT 8.36 1.95 9.51 2.12 ;
      RECT 9.18 2.12 9.51 2.98 ;
      RECT 6.425 2.73 6.76 2.905 ;
      RECT 6.425 2.65 6.675 2.73 ;
      RECT 7.46 2.29 7.63 2.905 ;
      RECT 5.905 0.92 6.235 1.09 ;
      RECT 5.905 0.75 9.025 0.92 ;
      RECT 8.775 0.92 9.965 1.09 ;
      RECT 5.905 0.6 6.235 0.75 ;
      RECT 6.905 0.35 7.155 0.75 ;
      RECT 7.835 0.35 8.085 0.75 ;
      RECT 8.775 0.35 9.025 0.75 ;
      RECT 9.715 0.35 9.965 0.92 ;
      RECT 2.395 0.35 6.235 0.6 ;
      RECT 3.335 0.6 3.505 0.84 ;
      RECT 0 3.245 10.08 3.415 ;
      RECT 8.73 2.29 8.98 3.245 ;
      RECT 9.71 1.95 9.96 3.245 ;
      RECT 0.115 1.95 0.365 3.245 ;
      RECT 1.065 2.29 1.395 3.245 ;
      RECT 3.025 2.73 3.355 3.245 ;
      RECT 2.025 2.39 2.355 3.245 ;
      RECT 5.925 2.39 6.255 3.245 ;
      RECT 6.405 0.085 6.735 0.58 ;
      RECT 0 -0.085 10.08 0.085 ;
      RECT 7.335 0.085 7.665 0.58 ;
      RECT 8.265 0.085 8.605 0.58 ;
      RECT 9.205 0.085 9.535 0.75 ;
    LAYER mcon ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
  END
END scs8ls_o221ai_4

MACRO scs8ls_o22a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.235 1.47 3.715 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 0.255 2.47 0.585 ;
        RECT 1.085 0.585 1.305 0.67 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B2

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.47 2.995 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.335 1.47 2.005 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.82 0.445 2.98 ;
        RECT 0.085 1.13 0.255 1.82 ;
        RECT 0.085 0.35 0.365 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.395 2.14 2.725 2.98 ;
      RECT 2.175 1.97 2.725 2.14 ;
      RECT 2.175 1.3 2.345 1.97 ;
      RECT 0.925 1.13 2.345 1.3 ;
      RECT 1.905 1.105 2.345 1.13 ;
      RECT 0.425 1.3 1.095 1.63 ;
      RECT 2.535 1.13 3.725 1.3 ;
      RECT 2.535 0.935 2.705 1.13 ;
      RECT 3.395 0.63 3.725 1.13 ;
      RECT 1.475 0.755 2.705 0.935 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 2.885 0.085 3.225 0.96 ;
      RECT 0.545 0.085 0.875 0.96 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 0.615 1.985 1.85 3.245 ;
      RECT 3.385 1.97 3.715 3.245 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_o22a_1

MACRO scs8ls_o22a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.3 3.735 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.71 1.43 3.235 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.43 1.875 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.43 2.5 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B2

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.82 0.865 1.13 ;
        RECT 0.635 1.13 0.805 1.82 ;
        RECT 0.535 0.35 0.79 0.82 ;
        RECT 0.635 1.82 0.965 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.465 0.96 3.725 1.13 ;
      RECT 2.465 0.52 2.795 0.96 ;
      RECT 3.475 0.35 3.725 0.96 ;
      RECT 1.505 0.35 2.795 0.52 ;
      RECT 1.505 0.52 1.835 0.71 ;
      RECT 2.35 2.12 2.68 2.94 ;
      RECT 1.135 1.95 2.68 2.12 ;
      RECT 1.135 0.88 2.295 1.13 ;
      RECT 2.005 0.8 2.295 0.88 ;
      RECT 1.135 1.63 1.305 1.95 ;
      RECT 0.975 1.3 1.305 1.63 ;
      RECT 1.135 1.13 1.305 1.3 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 0.965 0.085 1.295 0.64 ;
      RECT 2.965 0.085 3.295 0.79 ;
      RECT 0.105 0.085 0.365 1.13 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 1.135 2.29 1.79 3.245 ;
      RECT 3.4 1.95 3.73 3.245 ;
      RECT 0.135 1.82 0.465 3.245 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_o22a_2

MACRO scs8ls_nor2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.18 4.195 1.55 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 1.795 1.55 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.365 1.18 2.755 1.41 ;
        RECT 2.365 1.41 2.695 1.72 ;
        RECT 2.365 1.13 2.69 1.18 ;
        RECT 2.365 1.72 3.695 1.89 ;
        RECT 2.36 1.01 2.69 1.13 ;
        RECT 2.365 1.89 2.695 2.735 ;
        RECT 3.365 1.89 3.695 2.735 ;
        RECT 0.64 0.84 2.69 1.01 ;
        RECT 2.36 0.35 2.69 0.84 ;
        RECT 0.64 0.34 1.69 0.84 ;
    END
    ANTENNADIFFAREA 1.7936 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.915 2.905 4.145 3.075 ;
      RECT 3.865 1.82 4.145 2.905 ;
      RECT 1.915 1.89 2.195 2.905 ;
      RECT 0.115 1.72 2.195 1.89 ;
      RECT 0.115 1.89 0.445 2.98 ;
      RECT 1.015 1.89 1.345 2.98 ;
      RECT 2.865 2.06 3.195 2.905 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 0.645 2.06 0.815 3.245 ;
      RECT 1.545 2.06 1.715 3.245 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 2.86 0.085 4.205 1.01 ;
      RECT 0.115 0.085 0.47 1.01 ;
      RECT 1.86 0.085 2.19 0.67 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_nor2_4

MACRO scs8ls_nor2_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.415 1.65 5.695 1.78 ;
        RECT 4.415 1.78 4.745 2.735 ;
        RECT 5.365 1.78 5.695 2.735 ;
        RECT 4.415 1.48 7.545 1.65 ;
        RECT 6.265 1.65 6.595 2.735 ;
        RECT 7.215 1.65 7.545 2.735 ;
        RECT 4.415 1.31 6.275 1.48 ;
        RECT 4.26 1.18 6.275 1.31 ;
        RECT 1.86 1.14 6.275 1.18 ;
        RECT 1.86 1.01 5.275 1.14 ;
        RECT 5.945 0.35 6.275 1.14 ;
        RECT 1.86 0.35 2.19 1.01 ;
        RECT 3.26 0.35 3.59 1.01 ;
        RECT 4.26 0.35 5.275 1.01 ;
    END
    ANTENNADIFFAREA 2.8393 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.225 0.3 7.555 1.31 ;
    END
    ANTENNAGATEAREA 1.788 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.35 3.715 1.78 ;
    END
    ANTENNAGATEAREA 1.788 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 1.515 2.29 1.845 3.245 ;
      RECT 2.465 2.29 2.795 3.245 ;
      RECT 3.415 2.29 3.745 3.245 ;
      RECT 0.615 2.12 0.945 3.245 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 6.445 0.085 6.775 1.13 ;
      RECT 0.65 0.085 1.69 1.13 ;
      RECT 2.36 0.085 3.09 0.84 ;
      RECT 3.76 0.085 4.09 0.84 ;
      RECT 5.445 0.085 5.775 0.97 ;
      RECT 3.915 2.905 8.045 3.075 ;
      RECT 7.715 1.82 8.045 2.905 ;
      RECT 1.145 2.12 1.315 2.98 ;
      RECT 1.145 1.95 4.245 2.12 ;
      RECT 2.045 2.12 2.295 2.98 ;
      RECT 2.995 2.12 3.245 2.98 ;
      RECT 3.915 2.12 4.245 2.905 ;
      RECT 0.115 1.78 1.315 1.95 ;
      RECT 0.115 1.95 0.445 2.98 ;
      RECT 4.925 1.95 5.185 2.905 ;
      RECT 5.875 1.82 6.08 2.905 ;
      RECT 6.775 1.82 7.035 2.905 ;
    LAYER mcon ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_nor2_8

MACRO scs8ls_nor2b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035 1.18 1.365 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.875 1.82 2.315 2.98 ;
        RECT 2.145 1.15 2.315 1.82 ;
        RECT 1.535 0.98 2.315 1.15 ;
        RECT 1.535 0.35 1.785 0.98 ;
    END
    ANTENNADIFFAREA 0.6827 ;
  END Y

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.18 0.44 1.55 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END BN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.535 1.32 1.975 1.65 ;
      RECT 0.315 1.89 0.645 2.7 ;
      RECT 0.61 1.01 0.78 1.72 ;
      RECT 0.255 0.68 0.78 1.01 ;
      RECT 0.315 1.72 1.705 1.89 ;
      RECT 1.535 1.65 1.705 1.72 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 1.955 0.085 2.23 0.81 ;
      RECT 0.95 0.085 1.28 1.01 ;
      RECT 0 3.245 2.4 3.415 ;
      RECT 0.925 2.06 1.255 3.245 ;
    LAYER mcon ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nor2b_1

MACRO scs8ls_nor2b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.18 3.235 1.41 ;
        RECT 1.645 1.01 3.235 1.18 ;
        RECT 1.645 1.18 1.82 2.735 ;
        RECT 1.645 0.96 2.745 1.01 ;
        RECT 1.485 0.35 1.815 0.96 ;
        RECT 2.495 0.35 2.745 0.96 ;
    END
    ANTENNADIFFAREA 0.8244 ;
  END Y

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.53 1.47 0.86 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END BN

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.12 2.905 2.35 3.075 ;
      RECT 2.02 2.12 2.35 2.905 ;
      RECT 2.02 1.95 3.25 2.12 ;
      RECT 3 2.12 3.25 2.98 ;
      RECT 3 1.82 3.25 1.95 ;
      RECT 1.12 1.82 1.45 2.905 ;
      RECT 0.11 1.13 1.475 1.3 ;
      RECT 1.145 1.3 1.475 1.55 ;
      RECT 0.11 0.45 0.78 1.13 ;
      RECT 0.11 1.3 0.36 2.98 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.55 2.29 2.8 3.245 ;
      RECT 0.56 1.97 0.89 3.245 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.915 0.085 3.245 0.84 ;
      RECT 0.985 0.085 1.315 0.96 ;
      RECT 1.985 0.085 2.315 0.79 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_nor2b_2

MACRO scs8ls_nor2b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.84 0.355 1.41 ;
        RECT 0.185 1.41 0.355 1.51 ;
        RECT 0.125 0.67 3.81 0.84 ;
        RECT 0.185 1.51 0.705 1.58 ;
        RECT 2.06 0.53 2.39 0.67 ;
        RECT 3.56 0.51 3.81 0.67 ;
        RECT 0.185 1.58 2.055 1.68 ;
        RECT 0.535 1.68 2.055 1.75 ;
        RECT 1.885 1.75 2.055 1.85 ;
        RECT 1.885 1.85 2.165 2.06 ;
        RECT 1.885 2.06 3.145 2.23 ;
        RECT 1.885 2.23 2.165 2.735 ;
        RECT 2.895 2.23 3.145 2.735 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END Y

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.75 1.18 5.155 1.825 ;
    END
    ANTENNAGATEAREA 0.363 ;
  END BN

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.79 1.18 1.795 1.34 ;
        RECT 1.085 1.34 1.795 1.41 ;
        RECT 0.79 1.01 3.975 1.18 ;
        RECT 3.645 1.18 3.975 1.55 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.465 2.905 3.645 3.075 ;
      RECT 3.315 2.06 3.645 2.905 ;
      RECT 1.465 2.09 1.715 2.905 ;
      RECT 0.565 1.92 1.715 2.09 ;
      RECT 0.565 2.09 0.895 2.98 ;
      RECT 2.365 2.4 2.695 2.905 ;
      RECT 4.41 0.345 5.165 1.01 ;
      RECT 4.35 1.995 4.68 2.875 ;
      RECT 4.35 1.89 4.58 1.995 ;
      RECT 3.055 1.72 4.58 1.89 ;
      RECT 4.41 1.01 4.58 1.72 ;
      RECT 3.055 1.68 3.225 1.72 ;
      RECT 2.225 1.35 3.225 1.68 ;
      RECT 0 3.245 5.28 3.415 ;
      RECT 3.815 2.06 4.145 3.245 ;
      RECT 4.88 1.995 5.13 3.245 ;
      RECT 1.095 2.26 1.265 3.245 ;
      RECT 0.115 1.85 0.365 3.245 ;
      RECT 0 -0.085 5.28 0.085 ;
      RECT 3.99 0.085 4.24 0.84 ;
      RECT 1.55 0.085 1.88 0.5 ;
      RECT 2.57 0.085 3.38 0.5 ;
    LAYER mcon ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_nor2b_4

MACRO scs8ls_nor3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.36 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.87 1.3 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.3 1.815 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 2.12 1.815 2.98 ;
        RECT 0.53 1.95 1.815 2.12 ;
        RECT 0.53 1.13 0.7 1.95 ;
        RECT 0.53 0.88 1.805 1.13 ;
        RECT 0.615 0.365 0.805 0.88 ;
        RECT 1.475 0.35 1.805 0.88 ;
    END
    ANTENNADIFFAREA 0.7373 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.92 0.085 ;
      RECT 0.115 0.71 0.36 1.01 ;
      RECT 0.115 0.085 0.445 0.71 ;
      RECT 0.975 0.085 1.305 0.71 ;
      RECT 0 3.245 1.92 3.415 ;
      RECT 0.105 2.325 0.435 3.245 ;
      RECT 0.105 1.95 0.355 2.325 ;
    LAYER mcon ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nor3_1

MACRO scs8ls_nor3_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.18 0.975 1.55 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.18 3.255 1.38 ;
        RECT 1.305 1.38 3.255 1.55 ;
        RECT 1.305 1.22 1.635 1.38 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.65 0.31 3.235 0.98 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.35 0.445 0.84 ;
        RECT 0.115 0.84 1.98 1.01 ;
        RECT 0.115 1.01 0.355 1.72 ;
        RECT 1.65 1.01 1.98 1.05 ;
        RECT 1.65 0.35 1.98 0.84 ;
        RECT 0.115 1.72 0.945 1.89 ;
        RECT 0.615 1.89 0.945 2.735 ;
    END
    ANTENNADIFFAREA 0.8619 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.515 2.23 1.845 2.99 ;
      RECT 1.515 2.06 2.795 2.23 ;
      RECT 2.515 2.23 2.795 2.99 ;
      RECT 0.115 2.905 1.315 3.075 ;
      RECT 1.145 1.89 1.315 2.905 ;
      RECT 1.145 1.72 3.245 1.89 ;
      RECT 2.965 1.89 3.245 2.98 ;
      RECT 0.115 2.06 0.445 2.905 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.15 0.085 2.48 1.13 ;
      RECT 0.615 0.085 1.48 0.65 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.015 2.4 2.345 3.245 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_nor3_2

MACRO scs8ls_nor3_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 0.35 0.875 1.01 ;
        RECT 0.545 1.01 1.875 1.18 ;
        RECT 1.545 0.84 5.305 1.01 ;
        RECT 5.135 1.01 5.305 1.68 ;
        RECT 1.545 0.35 1.875 0.84 ;
        RECT 2.545 0.35 2.875 0.84 ;
        RECT 3.35 1.68 5.305 1.75 ;
        RECT 2.14 1.75 5.305 1.85 ;
        RECT 2.14 1.85 3.68 2 ;
    END
    ANTENNADIFFAREA 1.6748 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.785 0.34 5.635 0.67 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.18 4.965 1.35 ;
        RECT 1.31 1.35 4.965 1.51 ;
        RECT 1.31 1.51 2.755 1.52 ;
        RECT 1.31 1.52 1.64 1.68 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.92 1.795 2.17 ;
        RECT 1.625 2.17 6.135 2.19 ;
        RECT 0.605 1.35 0.935 1.92 ;
        RECT 1.625 2.19 4.02 2.34 ;
        RECT 3.85 2.02 6.135 2.17 ;
        RECT 5.805 0.33 6.135 2.02 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 6.72 3.415 ;
      RECT 5.835 2.7 6.165 3.245 ;
      RECT 0.56 2.68 0.89 3.245 ;
      RECT 0 -0.085 6.72 0.085 ;
      RECT 0.115 0.085 0.365 1.13 ;
      RECT 1.045 0.085 1.375 0.84 ;
      RECT 2.045 0.085 2.375 0.67 ;
      RECT 3.055 0.085 3.365 0.67 ;
      RECT 1.54 2.905 5.265 3.075 ;
      RECT 1.54 2.85 4.285 2.905 ;
      RECT 4.935 2.7 5.265 2.905 ;
      RECT 1.09 2.51 6.615 2.53 ;
      RECT 6.365 2.53 6.615 2.98 ;
      RECT 4.485 2.36 6.615 2.51 ;
      RECT 6.365 1.82 6.615 2.36 ;
      RECT 0.11 2.51 0.36 2.98 ;
      RECT 0.11 1.82 0.36 2.34 ;
      RECT 1.09 2.68 1.34 2.98 ;
      RECT 0.11 2.34 1.34 2.51 ;
      RECT 1.09 2.53 4.735 2.68 ;
      RECT 4.485 2.68 4.735 2.735 ;
      RECT 5.465 2.53 5.635 3 ;
    LAYER mcon ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_nor3_4

MACRO scs8ls_nor3b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.555 1.35 1.885 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985 1.35 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.18 0.815 1.55 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END CN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.33 0.35 2.795 1.01 ;
        RECT 1.33 1.01 2.795 1.18 ;
        RECT 2.625 1.18 2.795 2.29 ;
        RECT 1.33 0.35 1.66 1.01 ;
        RECT 2.275 2.29 2.795 2.98 ;
    END
    ANTENNADIFFAREA 0.7781 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.125 1.35 2.455 1.68 ;
      RECT 0.105 2.12 0.595 2.7 ;
      RECT 0.105 1.82 0.595 1.95 ;
      RECT 0.105 0.68 0.65 1.01 ;
      RECT 0.105 1.01 0.275 1.82 ;
      RECT 0.105 1.95 2.295 2.12 ;
      RECT 2.125 1.68 2.295 1.95 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 0.835 2.29 1.165 3.245 ;
      RECT 0 -0.085 2.88 0.085 ;
      RECT 0.83 0.085 1.16 1.01 ;
      RECT 1.83 0.085 2.16 0.84 ;
    LAYER mcon ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
  END
END scs8ls_nor3b_1

MACRO scs8ls_nor3b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.45 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END CN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.12 0.77 2.695 0.94 ;
        RECT 1.565 0.94 2.695 0.96 ;
        RECT 1.12 0.35 1.395 0.77 ;
        RECT 2.505 0.35 2.695 0.77 ;
        RECT 1.565 0.96 4.185 1.13 ;
        RECT 1.64 1.13 1.81 2.735 ;
        RECT 3.925 0.35 4.185 0.96 ;
    END
    ANTENNADIFFAREA 1.0057 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.605 1.35 3.275 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.35 4.675 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 3.46 2.29 3.79 3.245 ;
      RECT 4.425 1.95 4.69 3.245 ;
      RECT 0.56 1.95 0.89 3.245 ;
      RECT 2.46 2.12 2.79 2.735 ;
      RECT 2.46 1.95 4.24 2.12 ;
      RECT 3.99 2.12 4.24 2.98 ;
      RECT 1.11 2.905 3.24 3.075 ;
      RECT 2.97 2.29 3.24 2.905 ;
      RECT 2.01 1.82 2.29 2.905 ;
      RECT 1.11 1.82 1.44 2.905 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 4.355 0.085 4.685 1.13 ;
      RECT 0.62 0.085 0.95 0.94 ;
      RECT 1.565 0.085 2.335 0.6 ;
      RECT 2.865 0.085 3.755 0.77 ;
      RECT 0.085 1.11 1.335 1.28 ;
      RECT 1.005 1.28 1.335 1.55 ;
      RECT 0.085 0.35 0.45 1.11 ;
      RECT 0.085 1.95 0.36 2.98 ;
      RECT 0.085 1.28 0.255 1.95 ;
    LAYER mcon ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nor3b_2

MACRO scs8ls_nor3b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.765 1.18 7.095 1.55 ;
    END
    ANTENNAGATEAREA 0.363 ;
  END CN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.815 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.44 1.22 6.595 1.55 ;
        RECT 6.365 1.18 6.595 1.22 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.18 2.275 1.82 ;
        RECT 2.045 1.82 3.72 2.07 ;
        RECT 0.615 1.15 2.275 1.18 ;
        RECT 0.615 1.05 3.805 1.15 ;
        RECT 0.615 1.01 5.935 1.05 ;
        RECT 1.615 0.98 5.935 1.01 ;
        RECT 0.615 0.35 0.945 1.01 ;
        RECT 1.615 0.35 1.945 0.98 ;
        RECT 2.625 0.35 2.795 0.98 ;
        RECT 3.475 0.88 5.935 0.98 ;
        RECT 3.475 0.35 3.805 0.88 ;
        RECT 4.475 0.35 4.805 0.88 ;
        RECT 5.605 0.35 5.935 0.88 ;
    END
    ANTENNADIFFAREA 1.9855 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.525 2.24 5.1 2.41 ;
      RECT 4.93 2.41 5.1 2.99 ;
      RECT 4.795 2.23 5.1 2.24 ;
      RECT 4.795 2.06 6.08 2.23 ;
      RECT 5.81 2.23 6.08 2.99 ;
      RECT 1.525 2.41 1.855 2.735 ;
      RECT 1.525 2.12 1.87 2.24 ;
      RECT 0.615 1.95 1.87 2.12 ;
      RECT 0.615 2.12 0.945 2.735 ;
      RECT 6.785 1.89 7.055 2.7 ;
      RECT 3.89 1.72 7.565 1.89 ;
      RECT 7.395 1.01 7.565 1.72 ;
      RECT 6.605 0.35 7.565 1.01 ;
      RECT 3.89 1.65 4.195 1.72 ;
      RECT 2.58 1.32 4.195 1.65 ;
      RECT 0 3.245 7.68 3.415 ;
      RECT 4.4 2.58 4.73 3.245 ;
      RECT 5.3 2.4 5.63 3.245 ;
      RECT 6.25 2.06 6.58 3.245 ;
      RECT 7.235 2.06 7.565 3.245 ;
      RECT 0 -0.085 7.68 0.085 ;
      RECT 6.105 0.085 6.435 1.01 ;
      RECT 0.115 0.085 0.445 1.13 ;
      RECT 1.115 0.085 1.445 0.84 ;
      RECT 2.115 0.085 2.445 0.81 ;
      RECT 2.975 0.085 3.305 0.81 ;
      RECT 3.975 0.085 4.305 0.71 ;
      RECT 4.975 0.085 5.435 0.68 ;
      RECT 0.115 2.905 2.37 3.075 ;
      RECT 2.04 2.75 2.37 2.905 ;
      RECT 2.04 2.58 4.17 2.75 ;
      RECT 2.94 2.75 3.27 2.91 ;
      RECT 3.84 2.75 4.17 2.91 ;
      RECT 1.145 2.29 1.315 2.905 ;
      RECT 0.115 1.95 0.445 2.905 ;
    LAYER mcon ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_nor3b_4

MACRO scs8ls_nor4_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.54 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.975 1.35 1.315 2.89 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.35 1.875 2.15 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 2.445 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END D

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.265 1.95 2.785 2.98 ;
        RECT 2.615 1.18 2.785 1.95 ;
        RECT 0.78 1.01 2.785 1.18 ;
        RECT 0.78 0.35 1.04 1.01 ;
        RECT 1.81 0.35 2.14 1.01 ;
    END
    ANTENNADIFFAREA 0.7448 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.88 0.085 ;
      RECT 2.31 0.085 2.64 0.84 ;
      RECT 0.21 0.085 0.61 1.01 ;
      RECT 1.21 0.085 1.54 0.84 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 0.255 1.82 0.585 3.245 ;
    LAYER mcon ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nor4_1

MACRO scs8ls_nor4_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615 1.84 1.385 2.15 ;
        RECT 0.085 1.67 1.385 1.84 ;
        RECT 0.085 1 0.255 1.67 ;
        RECT 0.085 0.98 2.88 1 ;
        RECT 1.55 1 2.88 1.15 ;
        RECT 0.085 0.83 1.88 0.98 ;
        RECT 2.55 0.35 2.88 0.98 ;
        RECT 1.55 0.35 1.88 0.83 ;
    END
    ANTENNADIFFAREA 0.808 ;
  END Y

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.33 0.435 0.66 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END D

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885 0.28 4.215 1.71 ;
        RECT 2.455 1.71 4.215 1.88 ;
        RECT 2.455 1.65 2.625 1.71 ;
        RECT 2.285 1.32 2.625 1.65 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.095 1.18 3.715 1.54 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END A

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.65 1.795 2.15 ;
        RECT 1.565 1.5 2.075 1.65 ;
        RECT 0.425 1.32 2.075 1.5 ;
        RECT 0.425 1.17 0.7 1.32 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END C

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.565 2.66 1.835 2.98 ;
      RECT 2.035 2.05 4.205 2.22 ;
      RECT 3.94 2.22 4.205 2.98 ;
      RECT 0.115 2.32 2.285 2.49 ;
      RECT 2.035 2.49 2.285 2.98 ;
      RECT 2.035 2.22 2.285 2.32 ;
      RECT 2.035 1.82 2.285 2.05 ;
      RECT 0.115 2.49 0.365 3 ;
      RECT 0.115 2.01 0.445 2.32 ;
      RECT 2.475 2.56 2.805 3 ;
      RECT 2.475 2.39 3.755 2.56 ;
      RECT 3.505 2.56 3.755 3 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 2.975 2.73 3.305 3.245 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 3.05 0.085 3.38 1.01 ;
      RECT 0.605 0.085 1.38 0.6 ;
      RECT 2.05 0.085 2.38 0.81 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_nor4_2

MACRO scs8ls_nor4_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.35 1.875 1.78 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.435 1.35 3.785 1.78 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.35 6.595 1.78 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805 1.18 8.515 1.3 ;
        RECT 7.045 1.3 8.515 1.63 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.355 1.95 ;
        RECT 0.125 1.95 1.895 2.12 ;
        RECT 0.125 1.13 4.59 1.18 ;
        RECT 0.615 2.12 0.945 2.735 ;
        RECT 1.565 2.12 1.895 2.735 ;
        RECT 0.125 1.01 7.57 1.13 ;
        RECT 0.615 0.35 1.74 1.01 ;
        RECT 2.41 0.35 3.59 1.01 ;
        RECT 4.26 0.96 7.86 1.01 ;
        RECT 4.26 0.35 4.59 0.96 ;
        RECT 7.24 0.34 7.86 0.96 ;
    END
    ANTENNADIFFAREA 3.2144 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 6.695 2.29 7.025 3.245 ;
      RECT 7.695 2.29 8.025 3.245 ;
      RECT 4.375 2.12 4.625 2.735 ;
      RECT 4.375 1.95 8.525 2.12 ;
      RECT 5.34 2.12 5.56 2.735 ;
      RECT 6.255 2.12 6.525 2.98 ;
      RECT 7.195 2.12 7.525 2.98 ;
      RECT 8.195 2.12 8.525 2.98 ;
      RECT 8.195 1.82 8.525 1.95 ;
      RECT 2.465 2.905 6.075 3.075 ;
      RECT 4.825 2.3 5.155 2.905 ;
      RECT 5.745 2.3 6.075 2.905 ;
      RECT 2.465 2.29 2.795 2.905 ;
      RECT 3.365 2.29 3.695 2.905 ;
      RECT 0.115 2.905 2.265 3.075 ;
      RECT 2.095 2.12 2.265 2.905 ;
      RECT 2.095 1.95 4.145 2.12 ;
      RECT 2.97 2.12 3.19 2.735 ;
      RECT 3.895 2.12 4.145 2.735 ;
      RECT 2.095 1.82 2.265 1.95 ;
      RECT 0.115 2.29 0.445 2.905 ;
      RECT 1.145 2.29 1.395 2.905 ;
      RECT 0 -0.085 8.64 0.085 ;
      RECT 8.03 0.085 8.36 1.01 ;
      RECT 0.115 0.085 0.445 0.84 ;
      RECT 1.91 0.085 2.24 0.84 ;
      RECT 3.76 0.085 4.09 0.84 ;
      RECT 4.76 0.085 7.07 0.79 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
  END
END scs8ls_nor4_4

MACRO scs8ls_nor4b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 2.395 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.35 1.855 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985 1.35 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.11 0.815 1.44 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END DN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.85 3.275 2.98 ;
        RECT 3.105 1.18 3.275 1.85 ;
        RECT 1.29 1.01 3.275 1.18 ;
        RECT 1.29 0.35 1.62 1.01 ;
        RECT 2.3 0.35 2.63 1.01 ;
    END
    ANTENNADIFFAREA 0.8792 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.565 1.35 2.935 1.68 ;
      RECT 0.105 2.12 0.595 2.7 ;
      RECT 0.105 1.82 0.595 1.95 ;
      RECT 0.105 0.35 0.62 0.94 ;
      RECT 0.105 0.94 0.275 1.82 ;
      RECT 0.105 1.95 2.735 2.12 ;
      RECT 2.565 1.68 2.735 1.95 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 0.835 2.29 1.165 3.245 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.8 0.085 3.13 0.84 ;
      RECT 0.79 0.085 1.12 0.94 ;
      RECT 1.79 0.085 2.12 0.84 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_nor4b_1

MACRO scs8ls_nor4b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.44 0.35 3.77 1.01 ;
        RECT 2.44 1.01 5.145 1.18 ;
        RECT 2.925 1.18 3.095 1.95 ;
        RECT 2.44 0.96 2.77 1.01 ;
        RECT 4.815 0.35 5.145 1.01 ;
        RECT 1.655 1.95 3.095 2.12 ;
        RECT 1.25 0.79 2.77 0.96 ;
        RECT 1.655 2.12 1.825 2.735 ;
        RECT 1.655 1.82 1.825 1.95 ;
        RECT 2.44 0.35 2.77 0.79 ;
        RECT 1.25 0.33 1.58 0.79 ;
    END
    ANTENNADIFFAREA 1.3239 ;
  END Y

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 1.47 0.865 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END DN

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.295 1.35 4.195 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.35 5.635 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 4.835 2.29 5.165 3.245 ;
      RECT 0.565 1.97 0.895 3.245 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 5.315 0.085 5.645 1.13 ;
      RECT 0.75 0.085 1.08 0.96 ;
      RECT 1.75 0.085 2.27 0.6 ;
      RECT 2.94 0.085 3.27 0.84 ;
      RECT 3.94 0.085 4.645 0.79 ;
      RECT 2.025 2.29 3.255 2.46 ;
      RECT 3.005 2.46 3.255 2.735 ;
      RECT 1.125 1.82 1.455 2.905 ;
      RECT 1.125 2.905 2.275 3.075 ;
      RECT 2.025 2.46 2.275 2.905 ;
      RECT 2.475 2.905 4.265 3.075 ;
      RECT 2.475 2.63 2.805 2.905 ;
      RECT 3.935 2.29 4.265 2.905 ;
      RECT 3.485 2.12 3.735 2.735 ;
      RECT 3.485 1.95 5.625 2.12 ;
      RECT 4.465 2.12 4.635 2.98 ;
      RECT 5.375 2.12 5.625 2.98 ;
      RECT 0.115 1.13 1.775 1.3 ;
      RECT 1.105 1.3 1.775 1.55 ;
      RECT 0.115 0.35 0.58 1.13 ;
      RECT 0.115 1.3 0.365 2.98 ;
    LAYER mcon ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_nor4b_2

MACRO scs8ls_nor4b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405 1.18 5.635 1.95 ;
        RECT 2.025 1.95 5.635 1.99 ;
        RECT 3.5 1.01 9.465 1.18 ;
        RECT 2.025 1.99 2.355 2.735 ;
        RECT 2.975 1.99 5.635 2.12 ;
        RECT 2.025 1.82 3.305 1.95 ;
        RECT 3.5 1.18 3.75 1.3 ;
        RECT 3.5 0.35 3.75 1.01 ;
        RECT 4.905 0.35 5.235 1.01 ;
        RECT 6.25 0.35 6.58 1.01 ;
        RECT 7.25 0.35 7.58 1.01 ;
        RECT 8.275 0.35 8.525 1.01 ;
        RECT 9.215 0.35 9.465 1.01 ;
        RECT 2.975 2.12 3.305 2.735 ;
        RECT 2.5 1.3 3.75 1.47 ;
        RECT 2.5 1.15 2.83 1.3 ;
        RECT 1.57 0.98 2.83 1.15 ;
        RECT 1.57 0.35 1.82 0.98 ;
        RECT 2.5 0.35 2.83 0.98 ;
    END
    ANTENNADIFFAREA 2.4406 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805 1.35 9.475 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.35 7.555 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.92 1.35 5.155 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END C

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.92 0.55 1.93 ;
    END
    ANTENNAGATEAREA 0.363 ;
  END DN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 10.08 0.085 ;
      RECT 9.635 0.085 9.965 1.13 ;
      RECT 1.06 0.085 1.39 1.13 ;
      RECT 2 0.085 2.33 0.79 ;
      RECT 3 0.085 3.33 1.13 ;
      RECT 3.93 0.085 4.735 0.84 ;
      RECT 5.405 0.085 6.08 0.84 ;
      RECT 6.75 0.085 7.08 0.805 ;
      RECT 7.75 0.085 8.105 0.805 ;
      RECT 8.705 0.085 9.035 0.805 ;
      RECT 3.925 2.905 7.715 3.075 ;
      RECT 3.925 2.66 4.255 2.905 ;
      RECT 4.925 2.63 5.255 2.905 ;
      RECT 6.435 2.29 6.765 2.905 ;
      RECT 7.465 2.29 7.715 2.905 ;
      RECT 3.475 2.32 5.705 2.46 ;
      RECT 5.44 2.46 5.705 2.54 ;
      RECT 4.425 2.29 5.705 2.32 ;
      RECT 1.575 1.82 1.825 2.905 ;
      RECT 2.525 2.16 2.805 2.905 ;
      RECT 1.575 2.905 3.755 3.075 ;
      RECT 3.475 2.49 3.755 2.905 ;
      RECT 3.475 2.46 4.755 2.49 ;
      RECT 4.425 2.49 4.755 2.72 ;
      RECT 0.72 1.32 2.33 1.65 ;
      RECT 0.565 2.1 0.895 2.98 ;
      RECT 0.72 1.65 0.89 2.1 ;
      RECT 0.72 0.75 0.89 1.32 ;
      RECT 0.275 0.42 0.89 0.75 ;
      RECT 0 3.245 10.08 3.415 ;
      RECT 8.285 2.29 8.535 3.245 ;
      RECT 9.265 2.29 9.515 3.245 ;
      RECT 0.115 2.1 0.365 3.245 ;
      RECT 1.075 2.1 1.345 3.245 ;
      RECT 5.935 2.12 6.265 2.735 ;
      RECT 5.935 1.95 9.965 2.12 ;
      RECT 6.935 2.12 7.265 2.735 ;
      RECT 7.885 2.12 8.115 2.98 ;
      RECT 8.735 2.12 9.065 2.98 ;
      RECT 9.715 2.12 9.965 2.98 ;
      RECT 9.715 1.82 9.965 1.95 ;
    LAYER mcon ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nor4b_4

MACRO scs8ls_nor4bb_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.86 0.35 3.235 0.88 ;
        RECT 1.445 0.88 3.235 1.05 ;
        RECT 1.445 1.05 1.775 1.13 ;
        RECT 1.445 0.35 1.775 0.88 ;
        RECT 1.575 1.13 1.745 2.06 ;
        RECT 1.575 2.06 3.455 2.39 ;
    END
    ANTENNADIFFAREA 0.8484 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.075 1.35 1.405 2.15 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.915 1.35 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.435 1.55 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END CN

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.45 4.345 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END DN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 3.405 0.085 4.175 0.92 ;
      RECT 0.945 0.085 1.275 1.13 ;
      RECT 1.945 0.085 2.69 0.68 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 3.965 2.1 4.185 3.245 ;
      RECT 0.65 2.9 1.345 3.245 ;
      RECT 0.115 2.56 3.795 2.73 ;
      RECT 3.625 1.89 3.795 2.56 ;
      RECT 2.485 1.72 3.795 1.89 ;
      RECT 2.485 1.35 2.815 1.72 ;
      RECT 0.115 1.82 0.775 2.56 ;
      RECT 0.605 1.01 0.775 1.82 ;
      RECT 0.115 0.68 0.775 1.01 ;
      RECT 4.355 2.1 4.685 2.98 ;
      RECT 4.515 1.26 4.685 2.1 ;
      RECT 3.07 1.22 4.685 1.26 ;
      RECT 3.57 1.09 4.685 1.22 ;
      RECT 4.355 0.54 4.685 1.09 ;
      RECT 3.07 1.26 3.74 1.55 ;
    LAYER mcon ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
  END
END scs8ls_nor4bb_1

MACRO scs8ls_nor4bb_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.115 1.55 4.675 1.78 ;
        RECT 4.115 1.78 4.285 1.85 ;
        RECT 4.115 1.18 4.285 1.55 ;
        RECT 2.975 1.85 4.285 2.02 ;
        RECT 3.955 1.01 6.575 1.18 ;
        RECT 2.975 2.02 3.225 2.735 ;
        RECT 3.955 0.84 4.285 1.01 ;
        RECT 4.965 0.35 5.215 1.01 ;
        RECT 6.325 0.35 6.575 1.01 ;
        RECT 2.89 0.67 4.285 0.84 ;
        RECT 2.89 0.35 3.22 0.67 ;
        RECT 3.955 0.35 4.285 0.67 ;
    END
    ANTENNADIFFAREA 1.1981 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.86 1.35 6.115 1.635 ;
        RECT 5.405 1.635 6.115 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.31 1.35 7.075 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495 1.47 1.825 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END DN

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.47 1.315 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END CN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.495 1.01 3.785 1.18 ;
      RECT 3.615 1.18 3.785 1.35 ;
      RECT 3.615 1.35 3.945 1.68 ;
      RECT 0.485 0.71 2.665 0.88 ;
      RECT 2.495 0.88 2.665 1.01 ;
      RECT 0.115 1.13 0.815 1.3 ;
      RECT 0.485 0.88 0.815 1.13 ;
      RECT 0.485 0.36 0.815 0.71 ;
      RECT 0.115 1.97 0.445 2.98 ;
      RECT 0.115 1.3 0.285 1.97 ;
      RECT 2.155 1.35 3.165 1.68 ;
      RECT 1.885 2.14 2.215 2.98 ;
      RECT 1.885 1.97 2.325 2.14 ;
      RECT 2.155 1.68 2.325 1.97 ;
      RECT 2.155 1.3 2.325 1.35 ;
      RECT 1.62 1.05 2.325 1.3 ;
      RECT 2.495 2.905 3.725 3.075 ;
      RECT 3.395 2.36 3.725 2.905 ;
      RECT 3.395 2.19 4.675 2.36 ;
      RECT 4.345 2.36 4.675 2.735 ;
      RECT 2.495 1.85 2.775 2.905 ;
      RECT 3.895 2.905 5.685 3.075 ;
      RECT 3.895 2.53 4.175 2.905 ;
      RECT 5.355 2.29 5.685 2.905 ;
      RECT 4.905 2.12 5.155 2.735 ;
      RECT 4.905 1.95 7.085 2.12 ;
      RECT 5.855 2.12 6.185 2.98 ;
      RECT 6.755 2.12 7.085 2.98 ;
      RECT 4.905 1.82 5.155 1.95 ;
      RECT 0 3.245 7.2 3.415 ;
      RECT 6.385 2.29 6.555 3.245 ;
      RECT 0.615 1.97 1.715 3.245 ;
      RECT 0 -0.085 7.2 0.085 ;
      RECT 6.755 0.085 7.085 1.13 ;
      RECT 0.99 0.085 1.515 0.54 ;
      RECT 2.195 0.085 2.71 0.54 ;
      RECT 3.4 0.085 3.775 0.5 ;
      RECT 4.455 0.085 4.785 0.84 ;
      RECT 5.385 0.085 6.155 0.84 ;
    LAYER mcon ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_nor4bb_2

MACRO scs8ls_nor4bb_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 11.04 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN DN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.125 1.45 10.455 1.78 ;
    END
    ANTENNAGATEAREA 0.363 ;
  END DN

  PIN CN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.095 1.53 9.955 1.86 ;
    END
    ANTENNAGATEAREA 0.363 ;
  END CN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.705 0.35 8.035 0.885 ;
        RECT 6.445 0.885 8.035 1.055 ;
        RECT 6.445 1.055 6.615 1.3 ;
        RECT 6.445 0.35 6.775 0.885 ;
        RECT 5.525 1.3 6.615 1.47 ;
        RECT 5.99 1.47 6.32 1.725 ;
        RECT 5.525 1.085 5.775 1.3 ;
        RECT 5.99 1.725 7.23 2.055 ;
        RECT 2.665 1.01 5.775 1.085 ;
        RECT 0.615 0.915 5.775 1.01 ;
        RECT 0.615 1.01 0.945 1.13 ;
        RECT 0.615 0.84 2.915 0.915 ;
        RECT 3.595 0.35 3.845 0.915 ;
        RECT 4.515 0.35 4.845 0.915 ;
        RECT 5.525 0.35 5.775 0.915 ;
        RECT 0.615 0.35 0.945 0.84 ;
        RECT 1.615 0.35 1.945 0.84 ;
        RECT 2.665 0.35 2.915 0.84 ;
    END
    ANTENNADIFFAREA 2.5442 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.65 1.315 1.71 ;
        RECT 1.085 1.71 2.89 1.88 ;
        RECT 0.265 1.32 1.315 1.65 ;
        RECT 2.72 1.585 2.89 1.71 ;
        RECT 2.72 1.255 3.92 1.585 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.18 2.495 1.54 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.04 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.04 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 11.04 3.415 ;
      RECT 1.115 2.73 1.445 3.245 ;
      RECT 2.065 2.73 2.435 3.245 ;
      RECT 8.79 2.37 9.12 3.245 ;
      RECT 10.595 2.29 10.925 3.245 ;
      RECT 9.775 2.1 9.945 3.245 ;
      RECT 8.705 2.03 9.575 2.2 ;
      RECT 8.545 1.19 9.585 1.36 ;
      RECT 9.3 2.2 9.575 2.98 ;
      RECT 9.26 0.67 9.585 1.19 ;
      RECT 7.4 1.725 8.875 1.895 ;
      RECT 8.705 1.895 8.875 2.03 ;
      RECT 8.545 1.36 8.875 1.725 ;
      RECT 5.185 1.585 5.355 2.225 ;
      RECT 4.345 1.255 5.355 1.585 ;
      RECT 5.185 2.225 7.57 2.395 ;
      RECT 7.4 1.895 7.57 2.225 ;
      RECT 4.09 2.905 8.49 3.075 ;
      RECT 8.205 2.065 8.49 2.905 ;
      RECT 4.09 1.925 4.26 2.905 ;
      RECT 3.06 1.755 4.26 1.925 ;
      RECT 3.06 1.925 3.39 2.05 ;
      RECT 0.115 2.05 3.39 2.22 ;
      RECT 3.06 2.22 3.39 2.735 ;
      RECT 0.115 2.22 0.445 2.98 ;
      RECT 0.115 1.82 0.445 2.05 ;
      RECT 0 -0.085 11.04 0.085 ;
      RECT 8.205 0.085 8.75 0.68 ;
      RECT 10.095 0.085 10.495 0.94 ;
      RECT 0.115 0.085 0.445 1.13 ;
      RECT 1.115 0.085 1.445 0.67 ;
      RECT 2.115 0.085 2.445 0.67 ;
      RECT 3.085 0.085 3.415 0.745 ;
      RECT 4.015 0.085 4.345 0.745 ;
      RECT 5.015 0.085 5.345 0.745 ;
      RECT 5.945 0.085 6.275 1.13 ;
      RECT 6.945 0.085 7.535 0.68 ;
      RECT 4.47 2.565 8.035 2.735 ;
      RECT 7.76 2.065 8.035 2.565 ;
      RECT 4.47 1.755 4.8 2.565 ;
      RECT 0.615 2.56 0.945 2.98 ;
      RECT 0.615 2.39 2.885 2.56 ;
      RECT 1.645 2.56 1.895 2.98 ;
      RECT 2.635 2.56 2.885 2.905 ;
      RECT 2.635 2.905 3.89 3.075 ;
      RECT 3.56 2.095 3.89 2.905 ;
      RECT 10.145 2.12 10.395 2.98 ;
      RECT 10.145 1.95 10.925 2.12 ;
      RECT 10.755 1.28 10.925 1.95 ;
      RECT 9.755 1.11 10.925 1.28 ;
      RECT 10.665 0.35 10.925 1.11 ;
      RECT 9.755 0.425 9.925 1.11 ;
      RECT 8.92 0.255 9.925 0.425 ;
      RECT 8.92 0.425 9.09 0.85 ;
      RECT 8.205 0.85 9.09 1.02 ;
      RECT 8.205 1.02 8.375 1.225 ;
      RECT 6.785 1.225 8.375 1.555 ;
    LAYER mcon ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
  END
END scs8ls_nor4bb_4

MACRO scs8ls_o2111a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.82 0.445 2.98 ;
        RECT 0.095 1.04 0.265 1.82 ;
        RECT 0.095 0.35 0.355 1.04 ;
    END
    ANTENNADIFFAREA 0.5339 ;
  END X

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.55 1.335 1.88 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END D1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545 0.44 1.875 1.9 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END C1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.415 2.505 1.78 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END B1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.715 1.415 3.235 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.3 3.735 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.38 0.96 3.71 1.13 ;
      RECT 2.38 0.35 2.71 0.96 ;
      RECT 3.38 0.35 3.71 0.96 ;
      RECT 1.195 2.24 2.865 2.245 ;
      RECT 2.535 2.245 2.865 2.925 ;
      RECT 0.615 2.07 2.865 2.24 ;
      RECT 2.535 2.045 2.865 2.07 ;
      RECT 1.195 2.245 1.525 2.925 ;
      RECT 0.435 1.21 1.33 1.38 ;
      RECT 1.08 0.35 1.33 1.21 ;
      RECT 0.615 1.55 0.785 2.07 ;
      RECT 0.435 1.38 0.785 1.55 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 1.74 2.455 2.29 3.245 ;
      RECT 0.615 2.41 0.945 3.245 ;
      RECT 3.405 1.95 3.735 3.245 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 2.88 0.085 3.21 0.79 ;
      RECT 0.535 0.085 0.865 1.04 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o2111a_1

MACRO scs8ls_o2111a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.91 0.35 4.24 1.13 ;
        RECT 4.015 1.13 4.185 1.82 ;
        RECT 3.855 1.82 4.185 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.35 3.255 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END D1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.155 1.35 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END C1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.18 1.915 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.18 1.345 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.835 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.25 0.84 1.72 1.01 ;
      RECT 0.25 0.35 0.58 0.84 ;
      RECT 1.39 0.35 1.72 0.84 ;
      RECT 1.285 1.95 3.685 2.12 ;
      RECT 3.515 1.63 3.685 1.95 ;
      RECT 3.515 1.3 3.845 1.63 ;
      RECT 3.515 1.18 3.685 1.3 ;
      RECT 2.85 1.01 3.685 1.18 ;
      RECT 2.85 0.35 3.18 1.01 ;
      RECT 2.375 2.12 2.705 2.88 ;
      RECT 1.285 2.12 1.615 2.86 ;
      RECT 1.285 1.82 1.615 1.95 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 4.355 1.82 4.685 3.245 ;
      RECT 1.785 2.29 2.115 3.245 ;
      RECT 2.875 2.29 3.685 3.245 ;
      RECT 0.295 1.82 0.625 3.245 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 4.42 0.085 4.685 1.13 ;
      RECT 0.75 0.085 1.22 0.67 ;
      RECT 3.41 0.085 3.74 0.825 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o2111a_2

MACRO scs8ls_o2111a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805 1.18 8.035 1.48 ;
        RECT 7.295 1.48 8.035 1.65 ;
        RECT 6.185 1.01 8.035 1.18 ;
        RECT 7.295 1.65 7.545 1.85 ;
        RECT 6.185 0.35 6.515 1.01 ;
        RECT 7.185 0.35 7.515 1.01 ;
        RECT 6.315 1.85 7.545 2.18 ;
        RECT 6.315 2.18 6.59 2.98 ;
        RECT 7.295 2.18 7.545 2.98 ;
    END
    ANTENNADIFFAREA 1.1424 ;
  END X

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.325 1.45 5.655 1.78 ;
    END
    ANTENNAGATEAREA 0.522 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.45 5.155 1.78 ;
    END
    ANTENNAGATEAREA 0.522 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985 1.45 3.315 1.78 ;
    END
    ANTENNAGATEAREA 0.474 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.45 1.795 1.78 ;
    END
    ANTENNAGATEAREA 0.474 ;
  END C1

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.45 0.55 1.78 ;
    END
    ANTENNAGATEAREA 0.474 ;
  END D1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.365 1.28 2.775 1.3 ;
      RECT 2.365 1.11 5.505 1.28 ;
      RECT 2.365 1.05 3.555 1.11 ;
      RECT 4.235 0.52 4.565 1.11 ;
      RECT 5.335 0.35 5.505 1.11 ;
      RECT 3.305 0.52 3.555 1.05 ;
      RECT 1.41 0.88 1.74 1.13 ;
      RECT 1.41 0.71 3.125 0.88 ;
      RECT 1.41 0.595 1.74 0.71 ;
      RECT 2.875 0.52 3.125 0.71 ;
      RECT 0.115 0.6 0.38 1.115 ;
      RECT 0.115 0.425 1.23 0.6 ;
      RECT 1.06 0.6 1.23 1.13 ;
      RECT 0.115 0.255 2.25 0.425 ;
      RECT 1.92 0.425 2.25 0.54 ;
      RECT 3.72 2.46 4.05 2.735 ;
      RECT 3.72 2.29 5.61 2.46 ;
      RECT 5.28 2.46 5.61 2.98 ;
      RECT 5.975 1.35 7.125 1.68 ;
      RECT 0.115 1.95 6.145 2.12 ;
      RECT 5.975 1.68 6.145 1.95 ;
      RECT 3.22 2.905 4.55 3.075 ;
      RECT 4.22 2.63 4.55 2.905 ;
      RECT 3.22 2.12 3.55 2.905 ;
      RECT 1.115 2.12 1.445 2.82 ;
      RECT 2.15 2.12 2.48 2.82 ;
      RECT 2.15 1.94 2.48 1.95 ;
      RECT 0.115 2.12 0.445 2.82 ;
      RECT 0.72 1.13 0.89 1.95 ;
      RECT 0.55 0.77 0.89 1.13 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 7.685 0.085 8.015 0.815 ;
      RECT 3.735 0.085 4.065 0.94 ;
      RECT 4.825 0.085 5.155 0.94 ;
      RECT 5.685 0.085 6.015 1.13 ;
      RECT 6.685 0.085 7.015 0.815 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 7.715 1.82 8.045 3.245 ;
      RECT 4.78 2.63 5.11 3.245 ;
      RECT 0.615 2.315 0.945 3.245 ;
      RECT 1.615 2.315 1.945 3.245 ;
      RECT 2.685 2.315 3.015 3.245 ;
      RECT 5.815 2.29 6.145 3.245 ;
      RECT 6.765 2.35 7.095 3.245 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
  END
END scs8ls_o2111a_4

MACRO scs8ls_o2111ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.18 3.255 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.2 1.18 2.755 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.595 1.18 1.99 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 0.44 1.425 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END C1

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.58 1.18 0.91 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END D1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.88 1.89 1.315 2.98 ;
        RECT 0.115 1.72 2.315 1.89 ;
        RECT 1.985 1.89 2.315 2.98 ;
        RECT 0.115 1.01 0.285 1.72 ;
        RECT 0.115 0.35 0.785 1.01 ;
    END
    ANTENNADIFFAREA 1.1625 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.825 0.84 3.245 1.01 ;
      RECT 1.825 0.35 2.155 0.84 ;
      RECT 2.915 0.35 3.245 0.84 ;
      RECT 2.325 0.085 2.745 0.6 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.89 1.82 3.22 3.245 ;
      RECT 0.38 2.06 0.71 3.245 ;
      RECT 1.485 2.06 1.815 3.245 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_o2111ai_1

MACRO scs8ls_o2111ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.18 0.935 1.8 ;
        RECT 0.605 1.8 1.885 1.95 ;
        RECT 0.69 1.13 0.935 1.18 ;
        RECT 0.605 1.95 4.245 1.97 ;
        RECT 0.69 0.595 0.94 1.13 ;
        RECT 1.555 1.97 4.245 2.12 ;
        RECT 0.605 1.97 0.935 2.98 ;
        RECT 1.555 2.12 1.885 2.98 ;
        RECT 2.455 2.12 2.785 2.98 ;
        RECT 3.915 2.12 4.245 2.735 ;
    END
    ANTENNADIFFAREA 1.5512 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.35 5.635 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.35 4.675 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.35 3.715 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.18 1.795 1.3 ;
        RECT 1.345 1.3 2.015 1.63 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END C1

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.435 1.55 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END D1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.12 1.01 1.29 1.13 ;
      RECT 1.12 0.84 2.3 1.01 ;
      RECT 1.97 1.01 2.3 1.13 ;
      RECT 1.97 0.595 2.3 0.84 ;
      RECT 1.12 0.425 1.29 0.84 ;
      RECT 0.18 0.255 1.29 0.425 ;
      RECT 0.18 0.425 0.51 1.01 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 4.815 2.29 5.145 3.245 ;
      RECT 0.155 1.82 0.405 3.245 ;
      RECT 1.105 2.14 1.355 3.245 ;
      RECT 2.085 2.29 2.255 3.245 ;
      RECT 2.985 2.29 3.235 3.245 ;
      RECT 3.89 0.085 4.22 0.84 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 4.84 0.085 5.17 0.84 ;
      RECT 3.465 2.905 4.615 3.075 ;
      RECT 4.445 2.12 4.615 2.905 ;
      RECT 4.445 1.95 5.645 2.12 ;
      RECT 5.315 2.12 5.645 2.98 ;
      RECT 3.465 2.29 3.715 2.905 ;
      RECT 2.53 1.01 5.6 1.18 ;
      RECT 2.53 0.595 2.86 1.01 ;
      RECT 3.54 0.35 3.71 1.01 ;
      RECT 4.42 0.35 4.67 1.01 ;
      RECT 5.35 0.35 5.6 1.01 ;
      RECT 1.47 0.425 1.8 0.67 ;
      RECT 1.47 0.255 3.36 0.425 ;
      RECT 3.03 0.425 3.36 0.84 ;
    LAYER mcon ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_o2111ai_2

MACRO scs8ls_o2111ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.35 1.78 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END D1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.63 4.195 1.78 ;
        RECT 2.21 1.3 4.195 1.63 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END C1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805 1.35 9.49 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.285 1.35 7.635 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.35 6.115 1.78 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.55 2.04 1.78 ;
        RECT 1.87 1.78 2.04 1.8 ;
        RECT 1.565 1.13 1.805 1.55 ;
        RECT 1.87 1.8 3.52 1.95 ;
        RECT 0.615 0.77 1.805 1.13 ;
        RECT 0.115 1.95 9.515 1.97 ;
        RECT 0.115 1.97 2.2 2.12 ;
        RECT 3.19 1.97 9.515 2.12 ;
        RECT 0.115 2.12 1.2 2.98 ;
        RECT 1.87 2.12 2.2 2.98 ;
        RECT 3.19 2.12 3.52 2.98 ;
        RECT 4.19 2.12 4.52 2.98 ;
        RECT 8.185 2.12 8.515 2.735 ;
        RECT 9.185 2.12 9.515 2.735 ;
    END
    ANTENNADIFFAREA 3.4118 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 5.475 0.645 5.805 0.68 ;
      RECT 2.335 0.35 5.805 0.645 ;
      RECT 1.985 0.815 3.955 1.13 ;
      RECT 1.985 0.6 2.155 0.815 ;
      RECT 0.115 0.35 2.155 0.6 ;
      RECT 0.115 0.6 0.445 1.13 ;
      RECT 5.045 1.13 9.965 1.18 ;
      RECT 4.185 1.01 9.965 1.13 ;
      RECT 4.185 0.85 6.305 1.01 ;
      RECT 6.985 0.35 7.155 1.01 ;
      RECT 7.845 0.35 8.095 1.01 ;
      RECT 8.775 0.35 9.025 1.01 ;
      RECT 9.715 0.35 9.965 1.01 ;
      RECT 4.185 0.815 4.515 0.85 ;
      RECT 5.975 0.35 6.305 0.85 ;
      RECT 7.685 2.905 9.965 3.075 ;
      RECT 9.715 1.82 9.965 2.905 ;
      RECT 4.75 2.46 6.165 2.98 ;
      RECT 4.75 2.29 8.015 2.46 ;
      RECT 6.785 2.46 7.115 2.98 ;
      RECT 7.685 2.46 8.015 2.905 ;
      RECT 8.685 2.29 9.015 2.905 ;
      RECT 0 3.245 10.08 3.415 ;
      RECT 1.37 2.29 1.7 3.245 ;
      RECT 2.37 2.14 3.02 3.245 ;
      RECT 3.69 2.29 4.02 3.245 ;
      RECT 6.335 2.63 6.585 3.245 ;
      RECT 7.315 2.63 7.485 3.245 ;
      RECT 6.475 0.085 6.805 0.82 ;
      RECT 0 -0.085 10.08 0.085 ;
      RECT 7.335 0.085 7.665 0.82 ;
      RECT 8.265 0.085 8.595 0.82 ;
      RECT 9.205 0.085 9.535 0.82 ;
    LAYER mcon ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
  END
END scs8ls_o2111ai_4

MACRO scs8ls_mux4_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.915 1.18 6.345 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.28 0.805 1.55 ;
        RECT 0.435 1.26 1.845 1.28 ;
        RECT 0.435 1.18 1.655 1.26 ;
        RECT 1.485 1.28 1.845 1.59 ;
        RECT 0.635 1.11 1.655 1.18 ;
        RECT 1.485 0.59 1.655 1.11 ;
        RECT 1.485 0.42 3.105 0.59 ;
        RECT 2.835 0.59 3.105 1.11 ;
        RECT 2.835 1.11 5.745 1.28 ;
        RECT 2.835 1.28 3.105 1.78 ;
        RECT 4.395 1.28 4.725 1.55 ;
        RECT 5.475 1.28 5.745 1.75 ;
    END
    ANTENNAGATEAREA 0.768 ;
  END S0

  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.9 1.45 7.555 1.78 ;
    END
    ANTENNAGATEAREA 0.507 ;
  END S1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.855 1.45 4.195 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A3

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.975 1.45 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315 1.45 3.685 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A0

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.65 0.44 9.98 1.82 ;
        RECT 9.65 1.82 10 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 0.095 2.105 0.385 2.15 ;
      RECT 0.095 1.965 5.185 2.105 ;
      RECT 2.015 2.105 2.305 2.15 ;
      RECT 4.895 2.105 5.185 2.15 ;
      RECT 0.095 1.92 0.385 1.965 ;
      RECT 2.015 1.92 2.305 1.965 ;
      RECT 4.895 1.92 5.185 1.965 ;
    LAYER li1 ;
      RECT 4.925 1.46 5.265 2.15 ;
      RECT 7.2 2.905 9.13 3.075 ;
      RECT 7.2 2.71 7.53 2.905 ;
      RECT 8.96 1.68 9.13 2.905 ;
      RECT 8.96 1.35 9.385 1.68 ;
      RECT 8.96 0.425 9.13 1.35 ;
      RECT 7.12 0.255 9.13 0.425 ;
      RECT 7.12 0.425 7.45 0.6 ;
      RECT 0.255 2.15 0.585 2.98 ;
      RECT 0.095 1.92 0.585 2.15 ;
      RECT 0.095 0.5 0.465 1.01 ;
      RECT 0.095 1.01 0.265 1.92 ;
      RECT 5.775 2.37 7.98 2.54 ;
      RECT 7.81 2.54 7.98 2.565 ;
      RECT 7.65 1.95 7.98 2.37 ;
      RECT 7.81 2.565 8.79 2.735 ;
      RECT 8.62 0.765 8.79 2.565 ;
      RECT 7.845 0.595 8.79 0.765 ;
      RECT 7.845 0.765 8.015 0.77 ;
      RECT 4.53 0.77 8.015 0.94 ;
      RECT 6.69 0.35 6.94 0.77 ;
      RECT 5.055 2.66 5.945 2.91 ;
      RECT 5.775 2.54 5.945 2.66 ;
      RECT 4.53 0.35 5.105 0.77 ;
      RECT 2.045 1.45 2.325 2.15 ;
      RECT 8.2 1.78 8.45 2.395 ;
      RECT 7.725 1.45 8.45 1.78 ;
      RECT 8.185 0.935 8.45 1.45 ;
      RECT 5.435 1.96 7.08 2.2 ;
      RECT 6.56 1.95 7.08 1.96 ;
      RECT 6.56 1.11 7.955 1.28 ;
      RECT 6.56 1.28 6.73 1.95 ;
      RECT 4.115 2.32 5.605 2.49 ;
      RECT 5.435 2.2 5.605 2.32 ;
      RECT 4.115 2.12 4.285 2.32 ;
      RECT 2.495 1.95 4.285 2.12 ;
      RECT 2.495 2.12 3.445 2.98 ;
      RECT 2.495 1.09 2.665 1.95 ;
      RECT 1.85 0.76 2.665 1.09 ;
      RECT 0 3.245 10.56 3.415 ;
      RECT 10.2 1.82 10.45 3.245 ;
      RECT 6.165 2.71 6.495 3.245 ;
      RECT 3.615 2.29 3.945 3.245 ;
      RECT 0.755 1.95 1.085 3.245 ;
      RECT 9.3 1.85 9.47 3.245 ;
      RECT 0 -0.085 10.56 0.085 ;
      RECT 10.16 0.085 10.41 1.26 ;
      RECT 6.14 0.085 6.47 0.6 ;
      RECT 9.3 0.085 9.47 1.18 ;
      RECT 3.445 0.085 3.925 0.94 ;
      RECT 0.82 0.085 1.15 0.94 ;
    LAYER mcon ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 4.955 1.95 5.125 2.12 ;
      RECT 0.155 1.95 0.325 2.12 ;
      RECT 2.075 1.95 2.245 2.12 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
  END
END scs8ls_mux4_2

MACRO scs8ls_mux4_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 16.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.445 1.13 16.675 1.8 ;
        RECT 14.875 1.8 16.675 1.97 ;
        RECT 15.065 0.96 16.675 1.13 ;
        RECT 14.875 1.97 15.205 2.98 ;
        RECT 15.825 1.97 16.155 2.98 ;
        RECT 15.065 0.35 15.315 0.96 ;
        RECT 15.925 0.35 16.175 0.96 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END X

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.295 1.435 8.515 1.775 ;
    END
    ANTENNAGATEAREA 1.263 ;
  END S0

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.725 1.445 10.435 1.775 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.765 1.26 9.475 1.775 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.45 0.89 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.47 2.355 1.8 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A0

  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.15 1.3 12.835 1.78 ;
        RECT 12.15 1.275 13.865 1.3 ;
        RECT 13.54 1.3 13.865 1.55 ;
        RECT 12.665 1.13 13.865 1.275 ;
    END
    ANTENNAGATEAREA 0.771 ;
  END S1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 16.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 16.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 1.95 4.645 2.12 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 1.95 11.845 2.12 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
    LAYER met1 ;
      RECT 4.415 2.105 4.705 2.15 ;
      RECT 4.415 1.965 11.905 2.105 ;
      RECT 11.615 2.105 11.905 2.15 ;
      RECT 4.415 1.92 4.705 1.965 ;
      RECT 11.615 1.92 11.905 1.965 ;
    LAYER li1 ;
      RECT 0.565 1.97 2.695 2.14 ;
      RECT 2.525 1.77 2.695 1.97 ;
      RECT 2.525 1.6 4.19 1.77 ;
      RECT 4.02 1.77 4.19 2.735 ;
      RECT 0.565 2.14 0.895 2.98 ;
      RECT 0.565 1.95 0.895 1.97 ;
      RECT 3.05 0.96 3.38 1.09 ;
      RECT 1.97 0.79 3.38 0.96 ;
      RECT 1.575 0.62 2.14 0.79 ;
      RECT 3.05 0.595 3.38 0.79 ;
      RECT 1.575 0.47 1.81 0.62 ;
      RECT 0.545 0.275 1.81 0.47 ;
      RECT 0.545 0.47 0.875 0.86 ;
      RECT 1.515 2.48 1.845 2.98 ;
      RECT 1.515 2.31 3.3 2.48 ;
      RECT 3.045 2.48 3.3 2.735 ;
      RECT 2.99 1.94 3.3 2.31 ;
      RECT 0 3.245 16.8 3.415 ;
      RECT 16.325 2.14 16.655 3.245 ;
      RECT 8.32 2.965 8.65 3.245 ;
      RECT 9.39 2.965 9.73 3.245 ;
      RECT 2.045 2.65 2.295 3.245 ;
      RECT 1.095 2.31 1.345 3.245 ;
      RECT 10.465 2.285 10.635 3.245 ;
      RECT 0.115 1.95 0.365 3.245 ;
      RECT 5.4 1.82 5.73 3.245 ;
      RECT 14.375 1.82 14.705 3.245 ;
      RECT 15.405 2.14 15.655 3.245 ;
      RECT 13.875 1.89 14.205 2.98 ;
      RECT 13.005 1.72 14.205 1.89 ;
      RECT 14.035 0.96 14.205 1.72 ;
      RECT 13.905 0.595 14.205 0.96 ;
      RECT 13.005 1.47 13.33 1.72 ;
      RECT 0 -0.085 16.8 0.085 ;
      RECT 16.355 0.085 16.685 0.79 ;
      RECT 14.715 0.085 14.885 1.13 ;
      RECT 15.495 0.085 15.745 0.79 ;
      RECT 8.495 0.085 8.825 0.41 ;
      RECT 9.435 0.085 9.685 0.75 ;
      RECT 10.295 0.085 10.545 1.03 ;
      RECT 0.115 1.03 1.37 1.28 ;
      RECT 1.045 0.64 1.37 1.03 ;
      RECT 0.115 0.085 0.365 1.03 ;
      RECT 1.98 0.085 2.31 0.45 ;
      RECT 5.375 0.085 5.705 1.13 ;
      RECT 11.645 0.935 13.175 0.96 ;
      RECT 12.325 0.79 13.175 0.935 ;
      RECT 12.86 0.595 13.175 0.79 ;
      RECT 11.645 1.105 11.975 2.395 ;
      RECT 11.645 0.96 12.495 1.105 ;
      RECT 10.805 2.905 12.975 3.075 ;
      RECT 12.645 2.4 12.975 2.905 ;
      RECT 10.805 2.115 10.975 2.905 ;
      RECT 6.94 2.035 10.975 2.115 ;
      RECT 5.96 1.945 10.975 2.035 ;
      RECT 10.715 0.425 10.885 1.945 ;
      RECT 10.715 0.255 11.815 0.425 ;
      RECT 6.875 0.595 7.985 0.765 ;
      RECT 7.735 0.765 7.985 0.925 ;
      RECT 6.94 2.115 7.125 2.735 ;
      RECT 5.96 2.035 6.21 2.905 ;
      RECT 5.96 1.865 7.125 1.945 ;
      RECT 6.94 1.265 7.125 1.865 ;
      RECT 6.875 1.195 7.125 1.265 ;
      RECT 5.935 1.025 7.125 1.195 ;
      RECT 6.875 0.765 7.125 1.025 ;
      RECT 5.935 0.585 6.185 1.025 ;
      RECT 6.41 2.905 8.15 3.075 ;
      RECT 7.98 2.795 8.15 2.905 ;
      RECT 6.41 2.205 6.74 2.905 ;
      RECT 7.98 2.625 10.265 2.795 ;
      RECT 9.935 2.795 10.265 2.98 ;
      RECT 9.935 2.285 10.265 2.625 ;
      RECT 8.155 0.92 10.115 1.09 ;
      RECT 9.865 0.35 10.115 0.92 ;
      RECT 7.305 1.095 8.325 1.265 ;
      RECT 8.155 1.09 8.325 1.095 ;
      RECT 7.305 0.935 7.555 1.095 ;
      RECT 14.375 1.3 16.21 1.63 ;
      RECT 11.985 0.255 14.545 0.425 ;
      RECT 13.345 0.425 13.675 0.96 ;
      RECT 14.375 0.425 14.545 1.3 ;
      RECT 11.145 1.03 11.475 2.565 ;
      RECT 11.055 0.765 11.475 1.03 ;
      RECT 11.145 2.565 12.475 2.735 ;
      RECT 12.145 2.23 12.475 2.565 ;
      RECT 12.145 1.95 12.475 2.06 ;
      RECT 11.055 0.62 12.155 0.765 ;
      RECT 12.145 2.06 13.475 2.23 ;
      RECT 13.145 2.23 13.475 2.98 ;
      RECT 11.055 0.595 12.675 0.62 ;
      RECT 11.985 0.425 12.675 0.595 ;
      RECT 6.365 0.425 6.695 0.855 ;
      RECT 6.365 0.255 8.325 0.425 ;
      RECT 8.155 0.425 8.325 0.58 ;
      RECT 8.155 0.58 9.255 0.75 ;
      RECT 9.005 0.35 9.255 0.58 ;
      RECT 7.31 2.455 7.64 2.735 ;
      RECT 7.31 2.285 9.185 2.455 ;
      RECT 4.95 1.68 5.2 2.98 ;
      RECT 4.715 1.535 5.2 1.68 ;
      RECT 4.715 1.365 6.705 1.535 ;
      RECT 6.035 1.535 6.705 1.695 ;
      RECT 4.715 1.35 5.2 1.365 ;
      RECT 4.945 0.35 5.2 1.35 ;
      RECT 2.525 2.905 4.72 3.075 ;
      RECT 2.525 2.65 2.86 2.905 ;
      RECT 3.49 1.94 3.82 2.905 ;
      RECT 4.375 1.92 4.72 2.905 ;
      RECT 4.375 1.18 4.545 1.92 ;
      RECT 4.375 0.425 4.715 1.18 ;
      RECT 2.54 0.255 4.715 0.425 ;
      RECT 2.54 0.425 2.87 0.62 ;
      RECT 3.605 0.425 3.775 1.09 ;
      RECT 2.525 1.3 4.205 1.43 ;
      RECT 1.55 1.26 4.205 1.3 ;
      RECT 1.55 1.13 2.695 1.26 ;
      RECT 3.955 0.595 4.205 1.26 ;
      RECT 1.55 0.96 1.8 1.13 ;
  END
END scs8ls_mux4_4

MACRO scs8ls_nand2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.18 1.335 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.18 0.835 2.98 ;
        RECT 0.665 1.01 0.835 1.18 ;
        RECT 0.665 0.84 1.28 1.01 ;
        RECT 0.95 0.35 1.28 0.84 ;
    END
    ANTENNADIFFAREA 0.5469 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.435 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 1.44 3.415 ;
      RECT 1.005 1.82 1.335 3.245 ;
      RECT 0.105 1.82 0.435 3.245 ;
      RECT 0 -0.085 1.44 0.085 ;
      RECT 0.13 0.085 0.46 1.01 ;
    LAYER mcon ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_nand2_1

MACRO scs8ls_nand2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.35 1.815 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.35 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.18 2.275 1.95 ;
        RECT 0.57 1.95 2.275 2.12 ;
        RECT 1.455 1.01 2.275 1.18 ;
        RECT 0.57 2.12 0.82 2.98 ;
        RECT 1.56 2.12 1.73 2.98 ;
        RECT 1.455 0.595 1.785 1.01 ;
    END
    ANTENNADIFFAREA 0.9162 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.105 0.255 2.285 0.425 ;
      RECT 1.955 0.425 2.285 0.84 ;
      RECT 0.115 1.01 1.275 1.18 ;
      RECT 1.105 0.425 1.275 1.01 ;
      RECT 0.115 0.35 0.365 1.01 ;
      RECT 0 3.245 2.4 3.415 ;
      RECT 1.93 2.29 2.26 3.245 ;
      RECT 0.12 1.82 0.37 3.245 ;
      RECT 1.02 2.29 1.35 3.245 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 0.545 0.085 0.875 0.84 ;
    LAYER mcon ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nand2_2

MACRO scs8ls_nand2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.35 3.795 1.78 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.51 1.35 2.275 1.68 ;
        RECT 1.085 1.68 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.18 4.195 1.95 ;
        RECT 0.615 1.95 4.195 2.12 ;
        RECT 2.335 1.01 4.195 1.18 ;
        RECT 0.615 2.12 1.66 2.98 ;
        RECT 2.33 2.12 3.705 2.98 ;
        RECT 2.335 0.61 2.665 1.01 ;
        RECT 3.335 0.61 3.705 1.01 ;
    END
    ANTENNADIFFAREA 3.2861 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.915 0.255 4.205 0.425 ;
      RECT 3.875 0.425 4.205 0.805 ;
      RECT 0.115 1.01 2.165 1.18 ;
      RECT 1.915 0.425 2.165 1.01 ;
      RECT 0.115 0.35 0.365 1.01 ;
      RECT 1.055 0.35 1.225 1.01 ;
      RECT 2.835 0.425 3.165 0.805 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 3.875 2.29 4.205 3.245 ;
      RECT 0.115 1.85 0.445 3.245 ;
      RECT 1.83 2.29 2.16 3.245 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 0.545 0.085 0.875 0.805 ;
      RECT 1.405 0.085 1.735 0.805 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_nand2_4

MACRO scs8ls_nand2_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.38 1.13 4.71 1.95 ;
        RECT 2.14 1.95 4.71 2.12 ;
        RECT 4.335 1.05 4.71 1.13 ;
        RECT 2.14 2.12 2.47 2.98 ;
        RECT 4.38 2.12 4.71 2.98 ;
        RECT 4.335 0.77 7.895 1.05 ;
        RECT 7.725 1.05 7.895 1.95 ;
        RECT 5.94 1.95 7.895 2.12 ;
        RECT 5.94 2.12 6.27 2.98 ;
        RECT 7.32 2.12 7.55 2.98 ;
    END
    ANTENNADIFFAREA 2.2848 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.965 1.55 7.555 1.78 ;
        RECT 5.185 1.22 7.555 1.55 ;
    END
    ANTENNAGATEAREA 1.56 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 4.195 1.78 ;
    END
    ANTENNAGATEAREA 1.56 ;
  END B

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.985 0.35 8.045 0.6 ;
      RECT 0.105 1.165 4.155 1.18 ;
      RECT 1.035 1.01 4.155 1.165 ;
      RECT 3.985 0.6 4.155 1.01 ;
      RECT 1.895 0.35 2.155 1.01 ;
      RECT 3.075 0.35 3.305 1.01 ;
      RECT 0.105 1.18 1.86 1.355 ;
      RECT 0.105 0.35 0.355 1.165 ;
      RECT 1.035 0.35 1.225 1.01 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 0.535 0.085 0.865 0.995 ;
      RECT 1.395 0.085 1.725 0.84 ;
      RECT 2.325 0.085 2.905 0.84 ;
      RECT 3.475 0.085 3.805 0.84 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 7.72 2.29 8.05 3.245 ;
      RECT 0.66 1.95 1.97 3.245 ;
      RECT 2.64 2.29 4.21 3.245 ;
      RECT 4.88 1.82 5.21 3.245 ;
      RECT 5.44 1.82 5.77 3.245 ;
      RECT 6.44 2.29 7.15 3.245 ;
    LAYER mcon ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nand2_8

MACRO scs8ls_nand2b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 2.29 2.255 2.46 ;
        RECT 1.085 2.46 1.565 2.98 ;
        RECT 2.085 1.13 2.255 2.29 ;
        RECT 1.855 0.35 2.255 1.13 ;
    END
    ANTENNADIFFAREA 0.7102 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.35 1.345 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.3 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END AN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.515 1.3 1.915 1.63 ;
      RECT 0.115 1.95 1.685 2.12 ;
      RECT 1.515 1.63 1.685 1.95 ;
      RECT 1.515 1.13 1.685 1.3 ;
      RECT 0.115 0.96 1.685 1.13 ;
      RECT 0.115 2.12 0.445 2.7 ;
      RECT 0.115 0.54 0.38 0.96 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 0.55 0.085 1.22 0.79 ;
      RECT 0 3.245 2.4 3.415 ;
      RECT 1.735 2.65 2.07 3.245 ;
      RECT 0.65 2.29 0.915 3.245 ;
    LAYER mcon ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nand2b_1

MACRO scs8ls_nand2b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 0.57 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END AN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.39 2.275 1.82 ;
        RECT 1.645 1.82 2.275 1.95 ;
        RECT 1.7 1.22 2.275 1.39 ;
        RECT 1.645 1.95 2.795 2.2 ;
        RECT 1.7 0.63 1.87 1.22 ;
    END
    ANTENNADIFFAREA 0.8792 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.35 2.775 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.305 2.37 3.245 2.54 ;
      RECT 3.075 1.13 3.245 2.37 ;
      RECT 2.915 0.35 3.245 1.13 ;
      RECT 1.19 0.255 2.38 0.425 ;
      RECT 2.05 0.425 2.38 1.05 ;
      RECT 1.305 0.97 1.475 2.37 ;
      RECT 1.19 0.425 1.52 0.97 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.56 0.085 2.73 1.13 ;
      RECT 0.615 0.085 0.875 0.84 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.015 2.71 2.345 3.245 ;
      RECT 2.915 2.71 3.245 3.245 ;
      RECT 0.725 2.29 1.095 3.245 ;
      RECT 0.115 2.12 0.445 2.86 ;
      RECT 0.115 1.95 0.975 2.12 ;
      RECT 0.805 1.47 0.975 1.95 ;
      RECT 0.805 1.18 1.135 1.47 ;
      RECT 0.115 1.14 1.135 1.18 ;
      RECT 0.115 1.01 0.975 1.14 ;
      RECT 0.115 0.35 0.445 1.01 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nand2b_2

MACRO scs8ls_nand2b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.63 5.655 1.78 ;
        RECT 3.845 1.3 5.655 1.63 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.265 1.95 5.145 2.15 ;
        RECT 2.265 1.85 4.195 1.95 ;
        RECT 2.265 2.15 2.875 2.98 ;
        RECT 4.815 2.15 5.145 2.98 ;
        RECT 3.285 1.26 3.655 1.85 ;
        RECT 1.625 1.09 3.655 1.26 ;
        RECT 1.625 0.635 1.885 1.09 ;
        RECT 2.555 0.635 2.88 1.09 ;
    END
    ANTENNADIFFAREA 1.6343 ;
  END Y

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.3 1.115 1.78 ;
    END
    ANTENNAGATEAREA 0.363 ;
  END AN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.98 0.96 5.645 1.13 ;
      RECT 3.98 0.92 4.31 0.96 ;
      RECT 5.315 0.35 5.645 0.96 ;
      RECT 3.05 0.75 4.31 0.92 ;
      RECT 3.05 0.425 3.38 0.75 ;
      RECT 4.05 0.33 4.31 0.75 ;
      RECT 1.195 0.255 3.38 0.425 ;
      RECT 1.195 0.425 1.455 0.79 ;
      RECT 2.055 0.425 2.385 0.92 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 5.315 1.95 5.6 3.245 ;
      RECT 0.435 1.95 1.06 3.245 ;
      RECT 1.765 1.85 2.095 3.245 ;
      RECT 3.045 2.32 4.645 3.245 ;
      RECT 1.285 1.43 3.075 1.68 ;
      RECT 1.23 1.95 1.56 2.7 ;
      RECT 1.285 1.68 1.455 1.95 ;
      RECT 1.285 1.13 1.455 1.43 ;
      RECT 0.135 0.96 1.455 1.13 ;
      RECT 0.135 0.35 0.385 0.96 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 3.55 0.085 3.88 0.58 ;
      RECT 4.48 0.085 5.145 0.79 ;
      RECT 0.565 0.085 0.895 0.79 ;
    LAYER mcon ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nand2b_4

MACRO scs8ls_nand3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.18 1.915 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015 0.44 1.345 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.89 1.045 2.98 ;
        RECT 0.605 1.72 2.255 1.89 ;
        RECT 1.735 1.89 2.255 2.98 ;
        RECT 2.085 1.01 2.255 1.72 ;
        RECT 1.71 0.84 2.255 1.01 ;
        RECT 1.71 0.35 2.04 0.84 ;
    END
    ANTENNADIFFAREA 0.8773 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.835 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END C

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 0.32 0.085 0.65 1.01 ;
      RECT 0 3.245 2.4 3.415 ;
      RECT 0.185 1.82 0.435 3.245 ;
      RECT 1.215 2.06 1.545 3.245 ;
    LAYER mcon ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nand3_1

MACRO scs8ls_nand3_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965 1.43 2.295 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.265 1.55 1.795 1.68 ;
        RECT 1.425 1.68 1.795 1.95 ;
        RECT 1.265 1.43 1.595 1.55 ;
        RECT 1.425 1.95 2.825 2.12 ;
        RECT 2.655 1.65 2.825 1.95 ;
        RECT 2.655 1.32 3.065 1.65 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.735 1.55 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565 2.29 2.795 2.46 ;
        RECT 1.515 2.46 1.845 2.98 ;
        RECT 0.565 2.46 0.895 2.98 ;
        RECT 2.525 2.46 2.795 2.98 ;
        RECT 0.565 1.82 1.095 2.29 ;
        RECT 0.925 1.26 1.095 1.82 ;
        RECT 0.925 1.09 2.275 1.26 ;
        RECT 1.945 0.935 2.275 1.09 ;
    END
    ANTENNADIFFAREA 1.2208 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.53 0.085 0.86 0.58 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.995 1.82 3.245 3.245 ;
      RECT 0.115 1.82 0.365 3.245 ;
      RECT 1.065 2.63 1.315 3.245 ;
      RECT 2.015 2.63 2.345 3.245 ;
      RECT 0.1 0.75 3.26 0.765 ;
      RECT 2.93 0.765 3.26 1.15 ;
      RECT 1.04 0.595 3.26 0.75 ;
      RECT 2.945 0.405 3.26 0.595 ;
      RECT 0.1 0.92 0.43 1.01 ;
      RECT 0.1 0.35 0.35 0.75 ;
      RECT 0.1 0.765 1.37 0.92 ;
      RECT 1.04 0.33 1.21 0.595 ;
      RECT 1.455 0.255 2.765 0.425 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nand3_2

MACRO scs8ls_nand3_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.355 1.95 ;
        RECT 0.125 1.95 4.29 2.12 ;
        RECT 0.125 1.01 1.725 1.18 ;
        RECT 0.615 2.12 1.365 2.98 ;
        RECT 2.035 2.12 2.365 2.98 ;
        RECT 3.96 2.12 4.29 2.98 ;
        RECT 2.035 1.82 2.365 1.95 ;
        RECT 3.96 1.82 4.29 1.95 ;
        RECT 0.535 0.595 0.865 1.01 ;
        RECT 1.395 0.595 1.725 1.01 ;
    END
    ANTENNADIFFAREA 2.0048 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.35 1.535 1.78 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.56 1.63 3.715 1.78 ;
        RECT 2.13 1.35 3.715 1.63 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.495 1.63 6.115 1.78 ;
        RECT 4.14 1.34 6.115 1.63 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END C

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 4.085 0.085 4.415 0.75 ;
      RECT 0 -0.085 6.24 0.085 ;
      RECT 4.945 0.085 5.275 0.75 ;
      RECT 5.805 0.085 6.135 1.17 ;
      RECT 0 3.245 6.24 3.415 ;
      RECT 4.46 1.95 5.765 3.245 ;
      RECT 0.115 2.29 0.445 3.245 ;
      RECT 1.535 2.29 1.865 3.245 ;
      RECT 2.535 2.29 3.79 3.245 ;
      RECT 2.255 0.92 5.625 1.17 ;
      RECT 2.255 0.595 2.585 0.92 ;
      RECT 3.115 0.595 3.445 0.92 ;
      RECT 4.585 0.39 4.775 0.92 ;
      RECT 5.455 0.39 5.625 0.92 ;
      RECT 0.105 0.255 3.875 0.425 ;
      RECT 1.905 0.425 2.075 1.17 ;
      RECT 2.755 0.425 2.945 0.75 ;
      RECT 3.615 0.425 3.875 0.75 ;
      RECT 0.105 0.425 0.355 0.84 ;
      RECT 1.045 0.425 1.215 0.84 ;
    LAYER mcon ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nand3_4

MACRO scs8ls_nand3b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.35 1.915 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.305 1.95 2.795 2.12 ;
        RECT 2.305 2.12 2.795 2.98 ;
        RECT 1.305 2.12 1.635 2.98 ;
        RECT 2.305 1.82 2.795 1.95 ;
        RECT 2.625 1.15 2.795 1.82 ;
        RECT 2.425 0.79 2.795 1.15 ;
        RECT 2.25 0.37 2.795 0.79 ;
    END
    ANTENNADIFFAREA 1.0068 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.35 1.345 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END C

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.35 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END AN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 0.805 1.95 1.135 3.245 ;
      RECT 1.805 2.29 2.135 3.245 ;
      RECT 0 -0.085 2.88 0.085 ;
      RECT 0.545 0.085 1.22 0.81 ;
      RECT 2.085 1.32 2.455 1.65 ;
      RECT 0.105 0.98 2.255 1.15 ;
      RECT 2.085 1.15 2.255 1.32 ;
      RECT 0.105 1.95 0.6 2.7 ;
      RECT 0.105 1.15 0.275 1.95 ;
      RECT 0.105 0.56 0.375 0.98 ;
    LAYER mcon ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nand3b_1

MACRO scs8ls_nand3b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.35 4.195 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.43 1.795 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END C

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.45 0.55 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END AN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.18 2.8 1.95 ;
        RECT 1.26 1.95 3.695 2.12 ;
        RECT 2.47 1.01 2.8 1.18 ;
        RECT 1.26 2.12 1.635 2.98 ;
        RECT 2.335 2.12 2.585 2.98 ;
        RECT 3.365 2.12 3.695 2.98 ;
    END
    ANTENNADIFFAREA 1.3328 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.53 0.085 0.82 0.91 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 1.435 0.085 1.765 0.58 ;
      RECT 3.96 0.5 4.22 1.18 ;
      RECT 1.975 0.33 4.22 0.5 ;
      RECT 2.025 1.35 2.355 1.68 ;
      RECT 0.305 2.12 0.635 2.98 ;
      RECT 0.305 1.95 0.89 2.12 ;
      RECT 0.72 1.26 0.89 1.95 ;
      RECT 0.1 0.45 0.35 1.09 ;
      RECT 0.1 1.09 2.195 1.26 ;
      RECT 2.025 1.26 2.195 1.35 ;
      RECT 1.005 0.75 3.79 0.84 ;
      RECT 2.97 0.84 3.79 1.18 ;
      RECT 1.935 0.67 3.79 0.75 ;
      RECT 1.005 0.84 2.105 0.92 ;
      RECT 1.005 0.33 1.255 0.75 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 3.875 1.95 4.205 3.245 ;
      RECT 0.83 2.29 1.075 3.245 ;
      RECT 1.805 2.29 2.135 3.245 ;
      RECT 2.79 2.29 3.12 3.245 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nand3b_2

MACRO scs8ls_nand3b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.13 0.8 5.345 1.13 ;
        RECT 4.925 1.13 5.155 1.82 ;
        RECT 4.925 0.77 5.345 0.8 ;
        RECT 3.75 1.82 5.85 1.95 ;
        RECT 2.685 1.95 5.85 2.14 ;
    END
    ANTENNADIFFAREA 1.8665 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.82 1.18 7.075 1.65 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.765 1.35 3.235 1.78 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END C

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.35 1.095 1.78 ;
    END
    ANTENNAGATEAREA 0.363 ;
  END AN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.615 2.31 6.23 2.48 ;
      RECT 6.06 1.99 6.23 2.31 ;
      RECT 6.06 1.82 7.415 1.99 ;
      RECT 7.245 1.01 7.415 1.82 ;
      RECT 5.945 0.84 7.415 1.01 ;
      RECT 0.085 0.58 1.79 0.67 ;
      RECT 1.46 0.39 1.79 0.58 ;
      RECT 0.085 0.67 2.97 0.75 ;
      RECT 1.46 0.75 2.97 0.84 ;
      RECT 2.64 0.39 2.97 0.67 ;
      RECT 0.615 2.12 0.785 2.31 ;
      RECT 0.085 1.95 0.785 2.12 ;
      RECT 0.085 0.75 0.255 1.95 ;
      RECT 3.6 1.3 4.61 1.63 ;
      RECT 0.425 1.01 3.77 1.18 ;
      RECT 3.6 1.18 3.77 1.3 ;
      RECT 0.955 1.95 1.435 2.14 ;
      RECT 1.265 1.18 1.435 1.95 ;
      RECT 0.425 0.92 0.755 1.01 ;
      RECT 0 -0.085 7.68 0.085 ;
      RECT 0.935 0.085 1.28 0.41 ;
      RECT 1.97 0.085 2.46 0.5 ;
      RECT 3.14 0.085 3.47 0.84 ;
      RECT 0 3.245 7.68 3.415 ;
      RECT 1.49 2.65 2.565 3.245 ;
      RECT 3.135 2.65 3.63 3.245 ;
      RECT 4.58 2.65 5.4 3.245 ;
      RECT 5.97 2.65 7.565 3.245 ;
      RECT 0.115 2.29 0.445 3.245 ;
      RECT 6.4 2.16 7.565 2.65 ;
      RECT 3.7 0.6 4.03 0.63 ;
      RECT 3.7 0.35 7.565 0.6 ;
      RECT 5.515 0.6 7.565 0.67 ;
    LAYER mcon ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nand3b_4

MACRO scs8ls_nand4_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.18 2.775 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.715 1.18 2.275 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575 1.18 0.905 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END D

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.875 1.89 2.265 2.15 ;
        RECT 0.875 2.15 1.205 2.98 ;
        RECT 1.935 2.15 2.265 2.98 ;
        RECT 0.235 1.82 2.265 1.89 ;
        RECT 0.235 1.72 1.205 1.82 ;
        RECT 0.235 1.01 0.405 1.72 ;
        RECT 0.235 0.84 2.74 1.01 ;
        RECT 2.41 0.35 2.74 0.84 ;
    END
    ANTENNADIFFAREA 0.9365 ;
  END Y

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.18 1.475 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END C

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.88 0.085 ;
      RECT 0.11 0.085 0.785 0.6 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 2.435 1.82 2.765 3.245 ;
      RECT 0.375 2.06 0.705 3.245 ;
      RECT 1.4 2.32 1.73 3.245 ;
    LAYER mcon ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nand4_1

MACRO scs8ls_nand4_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885 1.35 4.215 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.68 1.35 3.715 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.09 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.43 1.35 2.44 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.18 4.675 1.95 ;
        RECT 0.635 1.95 4.675 2.12 ;
        RECT 3.845 1.01 4.675 1.18 ;
        RECT 3.84 2.12 4.675 2.15 ;
        RECT 0.635 2.12 0.9 2.98 ;
        RECT 1.57 2.12 1.9 2.98 ;
        RECT 2.83 2.12 3.16 2.98 ;
        RECT 3.845 0.645 4.175 1.01 ;
        RECT 3.84 2.15 4.125 2.98 ;
    END
    ANTENNADIFFAREA 1.6332 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.555 0.255 4.675 0.425 ;
      RECT 4.345 0.425 4.675 0.84 ;
      RECT 2.555 0.425 2.815 0.84 ;
      RECT 3.485 0.425 3.675 1.13 ;
      RECT 1.495 1.01 3.315 1.18 ;
      RECT 2.985 0.645 3.315 1.01 ;
      RECT 1.495 0.595 1.825 1.01 ;
      RECT 0.115 1.01 1.315 1.18 ;
      RECT 1.145 0.425 1.315 1.01 ;
      RECT 0.115 0.35 0.445 1.01 ;
      RECT 1.145 0.255 2.325 0.425 ;
      RECT 1.995 0.425 2.325 0.84 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 0.615 0.085 0.945 0.84 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 4.295 2.32 4.625 3.245 ;
      RECT 0.115 1.95 0.45 3.245 ;
      RECT 1.07 2.29 1.4 3.245 ;
      RECT 2.08 2.29 2.65 3.245 ;
      RECT 3.33 2.29 3.66 3.245 ;
    LAYER mcon ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nand4_2

MACRO scs8ls_nand4_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.35 6.16 1.78 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END B

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285 1.13 8.515 1.95 ;
        RECT 1.82 1.95 8.515 2.12 ;
        RECT 6.745 0.88 8.515 1.13 ;
        RECT 1.82 2.12 2.15 2.98 ;
        RECT 2.82 2.12 3.43 2.98 ;
        RECT 4.67 2.12 5.28 2.98 ;
        RECT 7.32 2.12 8.01 2.98 ;
        RECT 6.815 0.8 7.005 0.88 ;
        RECT 7.755 0.8 7.945 0.88 ;
    END
    ANTENNADIFFAREA 3.3216 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.735 1.35 8.085 1.78 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END A

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.35 4.195 1.78 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END C

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 4.595 0.52 4.925 0.71 ;
      RECT 4.595 0.35 8.525 0.52 ;
      RECT 5.455 0.52 5.785 0.71 ;
      RECT 6.315 0.52 6.645 0.71 ;
      RECT 7.175 0.52 7.505 0.71 ;
      RECT 8.195 0.52 8.525 0.71 ;
      RECT 2.745 0.88 6.215 1.13 ;
      RECT 2.745 0.85 3.935 0.88 ;
      RECT 5.095 0.8 5.285 0.88 ;
      RECT 5.955 0.8 6.145 0.88 ;
      RECT 0 -0.085 8.64 0.085 ;
      RECT 0.615 0.085 0.945 0.84 ;
      RECT 1.615 0.085 1.945 0.84 ;
      RECT 0.115 1.01 2.575 1.18 ;
      RECT 2.245 0.68 2.575 1.01 ;
      RECT 0.115 0.35 0.445 1.01 ;
      RECT 1.115 0.35 1.445 1.01 ;
      RECT 2.245 0.35 4.365 0.68 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 8.19 2.29 8.52 3.245 ;
      RECT 0.115 1.95 1.65 3.245 ;
      RECT 2.32 2.29 2.65 3.245 ;
      RECT 3.6 2.29 4.5 3.245 ;
      RECT 5.45 2.29 7.14 3.245 ;
    LAYER mcon ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nand4_4

MACRO scs8ls_nand4b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.18 2.395 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.18 1.855 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.285 1.89 2.635 2.15 ;
        RECT 1.285 2.15 1.615 2.98 ;
        RECT 2.285 2.15 2.635 2.98 ;
        RECT 1.285 1.82 3.275 1.89 ;
        RECT 1.615 1.72 3.275 1.82 ;
        RECT 3.105 1.05 3.275 1.72 ;
        RECT 2.905 0.35 3.275 1.05 ;
    END
    ANTENNADIFFAREA 1.0124 ;
  END Y

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985 1.18 1.315 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END D

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.18 0.815 1.55 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END AN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.565 1.22 2.935 1.55 ;
      RECT 0.105 0.84 2.735 1.01 ;
      RECT 2.565 1.01 2.735 1.22 ;
      RECT 0.105 1.82 0.58 2.7 ;
      RECT 0.105 0.68 0.65 0.84 ;
      RECT 0.105 1.01 0.275 1.82 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 0.855 0.085 1.185 0.67 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.805 2.06 3.135 3.245 ;
      RECT 0.785 1.82 1.115 3.245 ;
      RECT 1.785 2.32 2.115 3.245 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nand4b_1

MACRO scs8ls_nand4b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 2.59 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.35 4.195 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.35 5.635 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END D

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.985 1.51 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END AN

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.18 3.235 1.82 ;
        RECT 2.76 1.82 3.235 1.95 ;
        RECT 1.535 1.01 3.235 1.18 ;
        RECT 1.55 1.95 5.19 2.12 ;
        RECT 1.535 0.8 1.895 1.01 ;
        RECT 1.55 2.12 1.825 2.98 ;
        RECT 2.76 2.12 3.09 2.98 ;
        RECT 3.76 2.12 4.09 2.98 ;
        RECT 4.86 2.12 5.19 2.98 ;
        RECT 1.55 1.85 1.825 1.95 ;
    END
    ANTENNADIFFAREA 1.5734 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.545 0.085 0.875 0.67 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 4.865 0.085 5.195 0.76 ;
      RECT 2.505 0.425 2.835 0.5 ;
      RECT 2.505 0.255 4.335 0.425 ;
      RECT 4.005 0.425 4.335 0.76 ;
      RECT 2.075 0.67 3.345 0.84 ;
      RECT 2.075 0.63 2.325 0.67 ;
      RECT 3.015 0.595 3.345 0.67 ;
      RECT 1.105 0.35 2.325 0.63 ;
      RECT 3.575 0.93 5.645 1.18 ;
      RECT 3.575 0.595 3.825 0.93 ;
      RECT 4.505 0.4 4.695 0.93 ;
      RECT 5.395 0.4 5.645 0.93 ;
      RECT 1.155 1.35 1.72 1.68 ;
      RECT 0.505 1.85 0.835 2.86 ;
      RECT 0.505 1.68 1.325 1.85 ;
      RECT 1.155 1.01 1.325 1.35 ;
      RECT 0.115 0.84 1.325 1.01 ;
      RECT 0.115 0.35 0.365 0.84 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 5.36 1.95 5.645 3.245 ;
      RECT 1.04 2.02 1.37 3.245 ;
      RECT 1.995 2.29 2.59 3.245 ;
      RECT 3.26 2.29 3.59 3.245 ;
      RECT 4.32 2.29 4.65 3.245 ;
    LAYER mcon ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nand4b_2

MACRO scs8ls_nand4b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805 1.3 9.015 1.78 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END D

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.26 4.675 1.82 ;
        RECT 2.395 1.13 4.675 1.26 ;
        RECT 4.31 1.82 4.675 1.95 ;
        RECT 1.535 1.09 4.675 1.13 ;
        RECT 2.05 1.95 8.505 2.12 ;
        RECT 1.535 0.88 2.725 1.09 ;
        RECT 2.05 2.12 2.67 2.98 ;
        RECT 4.37 2.12 4.59 2.98 ;
        RECT 6.065 2.12 6.66 2.98 ;
        RECT 8.215 2.12 8.505 2.98 ;
        RECT 2.05 1.85 2.68 1.95 ;
        RECT 2.395 0.595 2.725 0.88 ;
    END
    ANTENNADIFFAREA 2.6656 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.13 1.43 4.14 1.78 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.35 7.555 1.78 ;
    END
    ANTENNAGATEAREA 0.78 ;
  END C

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.3 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.363 ;
  END AN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.12 0.085 ;
      RECT 7.27 0.085 7.6 0.78 ;
      RECT 8.13 0.085 8.505 0.78 ;
      RECT 0.545 0.085 0.875 0.6 ;
      RECT 0 3.245 9.12 3.415 ;
      RECT 8.675 1.95 8.955 3.245 ;
      RECT 0.505 1.95 0.835 3.245 ;
      RECT 1.54 1.85 1.87 3.245 ;
      RECT 2.85 2.29 4.19 3.245 ;
      RECT 4.76 2.29 5.885 3.245 ;
      RECT 6.835 2.29 8.035 3.245 ;
      RECT 5.605 0.6 5.795 0.71 ;
      RECT 5.535 0.58 6.725 0.6 ;
      RECT 6.395 0.6 6.725 0.84 ;
      RECT 3.255 0.33 6.725 0.58 ;
      RECT 5.965 1.13 7.17 1.18 ;
      RECT 5.105 1.01 9.005 1.13 ;
      RECT 5.105 0.96 6.215 1.01 ;
      RECT 6.92 0.96 9.005 1.01 ;
      RECT 5.105 0.77 5.435 0.96 ;
      RECT 5.965 0.77 6.215 0.96 ;
      RECT 6.92 0.35 7.1 0.96 ;
      RECT 7.77 0.35 7.96 0.96 ;
      RECT 8.675 0.35 9.005 0.96 ;
      RECT 2.905 0.75 4.875 0.92 ;
      RECT 2.905 0.425 3.075 0.75 ;
      RECT 1.105 0.255 3.075 0.425 ;
      RECT 1.105 0.425 1.435 0.71 ;
      RECT 1.965 0.425 2.215 0.71 ;
      RECT 1.005 1.43 2.85 1.68 ;
      RECT 1.005 1.68 1.335 2.7 ;
      RECT 1.005 1.13 1.335 1.43 ;
      RECT 0.115 0.96 1.335 1.13 ;
      RECT 0.115 0.77 0.445 0.96 ;
    LAYER mcon ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
  END
END scs8ls_nand4b_4

MACRO scs8ls_nand4bb_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985 0.81 3.315 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.95 4.225 2.12 ;
        RECT 2.525 2.12 3.095 2.31 ;
        RECT 2.525 1.82 3.095 1.95 ;
        RECT 3.765 2.12 4.225 2.98 ;
        RECT 4.055 1.18 4.225 1.95 ;
        RECT 1.675 2.31 3.095 2.48 ;
        RECT 3.485 1.01 4.225 1.18 ;
        RECT 1.675 2.48 2.005 2.98 ;
        RECT 2.765 2.48 3.095 2.98 ;
        RECT 3.485 0.62 3.655 1.01 ;
        RECT 1.72 0.35 3.655 0.62 ;
    END
    ANTENNADIFFAREA 1.24865 ;
  END Y

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.35 3.885 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END D

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.255 0.48 0.67 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END AN

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.47 1.315 1.8 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END BN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.115 1.13 2.015 1.3 ;
      RECT 1.685 1.3 2.015 1.55 ;
      RECT 0.115 1.97 0.445 2.85 ;
      RECT 0.115 1.3 0.285 1.97 ;
      RECT 0.115 0.84 0.47 1.13 ;
      RECT 2.185 1.22 2.745 1.55 ;
      RECT 1.115 2.14 1.445 2.85 ;
      RECT 1.15 0.63 1.49 0.79 ;
      RECT 1.115 1.97 2.355 2.14 ;
      RECT 2.185 1.55 2.355 1.97 ;
      RECT 2.185 0.96 2.355 1.22 ;
      RECT 1.15 0.79 2.355 0.96 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 3.825 0.085 4.155 0.84 ;
      RECT 0.65 0.085 0.98 0.96 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 0.615 1.97 0.945 3.245 ;
      RECT 2.175 2.65 2.595 3.245 ;
      RECT 3.265 2.29 3.595 3.245 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_nand4bb_1

MACRO scs8ls_nand4bb_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.18 1.335 1.51 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END BN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.625 1.35 6.595 1.68 ;
        RECT 6.365 1.68 6.595 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.35 5.385 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END C

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.26 4.195 1.85 ;
        RECT 2.345 1.85 4.195 1.95 ;
        RECT 2.685 1.09 4.195 1.26 ;
        RECT 2.345 1.95 6.105 2.02 ;
        RECT 2.345 1.82 2.675 1.85 ;
        RECT 2.685 0.84 2.855 1.09 ;
        RECT 3.345 2.02 6.105 2.12 ;
        RECT 2.345 2.02 2.675 2.98 ;
        RECT 5.775 1.85 6.105 1.95 ;
        RECT 2.345 0.67 2.855 0.84 ;
        RECT 3.345 2.12 3.675 2.98 ;
        RECT 4.775 2.12 5.105 2.98 ;
        RECT 5.775 2.12 6.105 2.98 ;
    END
    ANTENNADIFFAREA 1.6145 ;
  END Y

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.3 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END AN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.345 1.43 3.795 1.6 ;
      RECT 3.125 1.6 3.795 1.68 ;
      RECT 1.185 1.82 1.675 2.07 ;
      RECT 1.505 1.18 1.675 1.82 ;
      RECT 1.13 0.35 1.675 1.01 ;
      RECT 1.505 1.01 2.515 1.18 ;
      RECT 2.345 1.18 2.515 1.43 ;
      RECT 0 3.245 6.72 3.415 ;
      RECT 6.275 1.95 6.605 3.245 ;
      RECT 0.65 2.58 0.98 3.245 ;
      RECT 1.845 2.58 2.175 3.245 ;
      RECT 2.845 2.19 3.175 3.245 ;
      RECT 3.845 2.29 4.605 3.245 ;
      RECT 5.275 2.29 5.605 3.245 ;
      RECT 0 -0.085 6.72 0.085 ;
      RECT 5.84 0.085 6.17 0.815 ;
      RECT 0.63 0.085 0.96 1.01 ;
      RECT 4.41 1.01 6.6 1.18 ;
      RECT 4.41 0.62 4.74 1.01 ;
      RECT 5.42 0.35 5.67 1.01 ;
      RECT 6.35 0.35 6.6 1.01 ;
      RECT 3.365 0.425 3.695 0.58 ;
      RECT 3.365 0.255 5.24 0.425 ;
      RECT 4.91 0.425 5.24 0.815 ;
      RECT 3.025 0.75 4.18 0.92 ;
      RECT 3.025 0.5 3.195 0.75 ;
      RECT 1.845 0.33 3.195 0.5 ;
      RECT 1.845 0.5 2.175 0.84 ;
      RECT 0.095 2.24 2.175 2.41 ;
      RECT 1.845 1.35 2.175 2.24 ;
      RECT 0.095 2.41 0.445 2.86 ;
      RECT 0.095 1.95 0.445 2.24 ;
      RECT 0.095 0.35 0.46 1.03 ;
      RECT 0.095 1.03 0.265 1.95 ;
    LAYER mcon ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_nand4bb_2

MACRO scs8ls_nand4bb_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 2.23 2.965 2.99 ;
        RECT 2.525 2.06 4.815 2.23 ;
        RECT 3.635 2.23 3.865 2.99 ;
        RECT 4.535 2.23 4.815 2.98 ;
        RECT 4.485 2.02 4.815 2.06 ;
        RECT 4.485 1.99 5.685 2.02 ;
        RECT 5.515 2.02 5.685 2.98 ;
        RECT 4.485 1.95 9.515 1.99 ;
        RECT 6.335 1.99 9.515 2.12 ;
        RECT 4.485 1.85 6.665 1.95 ;
        RECT 7.335 1.82 7.665 1.95 ;
        RECT 6.335 2.12 6.665 2.98 ;
        RECT 7.335 2.12 7.665 2.98 ;
        RECT 8.285 2.12 8.615 2.98 ;
        RECT 9.185 2.12 9.515 2.98 ;
        RECT 5.515 1.82 6.665 1.85 ;
        RECT 5.515 1.26 5.685 1.82 ;
        RECT 3.335 1.09 5.685 1.26 ;
        RECT 3.335 1.04 3.505 1.09 ;
        RECT 2.32 0.87 3.505 1.04 ;
        RECT 2.32 0.595 2.65 0.87 ;
        RECT 3.335 0.595 3.505 0.87 ;
    END
    ANTENNADIFFAREA 3.2361 ;
  END Y

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.55 1.795 1.88 ;
    END
    ANTENNAGATEAREA 0.363 ;
  END BN

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.44 1.45 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.363 ;
  END AN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.265 1.3 9.955 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845 1.65 7.075 1.78 ;
        RECT 6.185 1.32 7.61 1.65 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END C

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.685 0.75 5.895 0.92 ;
      RECT 5.565 0.595 5.895 0.75 ;
      RECT 3.685 0.425 3.935 0.75 ;
      RECT 1.93 0.255 3.935 0.425 ;
      RECT 1.93 0.425 2.1 1.04 ;
      RECT 2.82 0.425 3.15 0.7 ;
      RECT 4.115 0.425 5.385 0.58 ;
      RECT 4.115 0.255 7.745 0.425 ;
      RECT 6.555 0.425 6.885 0.81 ;
      RECT 7.415 0.425 7.745 0.81 ;
      RECT 1.59 1.21 3.165 1.38 ;
      RECT 2.155 1.38 3.165 1.55 ;
      RECT 0.1 0.66 1.76 0.83 ;
      RECT 1.59 0.83 1.76 1.21 ;
      RECT 0.645 2.12 0.815 2.98 ;
      RECT 0.1 1.95 0.815 2.12 ;
      RECT 0.1 0.83 0.445 1.28 ;
      RECT 0.1 0.55 0.445 0.66 ;
      RECT 0.1 1.28 0.27 1.95 ;
      RECT 6.125 1.13 8.095 1.15 ;
      RECT 6.125 0.98 9.965 1.13 ;
      RECT 6.125 0.595 6.375 0.98 ;
      RECT 7.065 0.595 7.235 0.98 ;
      RECT 7.925 0.96 9.965 0.98 ;
      RECT 7.925 0.35 8.095 0.96 ;
      RECT 8.785 0.35 8.955 0.96 ;
      RECT 9.635 0.35 9.965 0.96 ;
      RECT 4.145 1.43 5.345 1.68 ;
      RECT 1.515 2.22 1.795 2.98 ;
      RECT 1.125 2.05 2.135 2.22 ;
      RECT 1.965 1.89 2.135 2.05 ;
      RECT 1.965 1.72 4.315 1.89 ;
      RECT 4.145 1.68 4.315 1.72 ;
      RECT 1.125 1.33 1.295 2.05 ;
      RECT 1.125 1 1.42 1.33 ;
      RECT 0 3.245 10.08 3.415 ;
      RECT 9.715 1.95 9.965 3.245 ;
      RECT 1.015 2.39 1.345 3.245 ;
      RECT 2.005 2.39 2.335 3.245 ;
      RECT 0.115 2.29 0.445 3.245 ;
      RECT 3.135 2.4 3.465 3.245 ;
      RECT 4.035 2.4 4.365 3.245 ;
      RECT 4.985 2.19 5.315 3.245 ;
      RECT 5.885 2.16 6.135 3.245 ;
      RECT 6.835 2.29 7.165 3.245 ;
      RECT 7.865 2.29 8.115 3.245 ;
      RECT 8.815 2.29 8.985 3.245 ;
      RECT 0 -0.085 10.08 0.085 ;
      RECT 8.275 0.085 8.605 0.79 ;
      RECT 9.135 0.085 9.465 0.79 ;
      RECT 0.625 0.085 0.955 0.49 ;
    LAYER mcon ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
  END
END scs8ls_nand4bb_4

MACRO scs8ls_nor2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.3 0.455 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.645 1.95 1.315 2.89 ;
        RECT 0.985 2.89 1.315 2.98 ;
        RECT 0.645 1.13 0.815 1.95 ;
        RECT 0.565 0.35 0.815 1.13 ;
    END
    ANTENNADIFFAREA 0.5376 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985 1.3 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 1.44 3.415 ;
      RECT 0.115 1.95 0.445 3.245 ;
      RECT 0 -0.085 1.44 0.085 ;
      RECT 0.995 0.085 1.325 1.13 ;
      RECT 0.135 0.085 0.385 1.13 ;
    LAYER mcon ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_nor2_1

MACRO scs8ls_nor2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805 0.44 2.275 1.41 ;
        RECT 1.805 1.41 2.135 1.605 ;
        RECT 1.805 0.255 2.135 0.44 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.82 0.945 2.735 ;
        RECT 0.615 0.35 0.945 1.82 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END Y

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.18 0.445 1.55 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END B

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.155 2.905 1.305 3.075 ;
      RECT 1.135 1.945 1.305 2.905 ;
      RECT 1.135 1.775 2.285 1.945 ;
      RECT 1.955 1.945 2.285 2.98 ;
      RECT 0.155 1.82 0.405 2.905 ;
      RECT 0 3.245 2.4 3.415 ;
      RECT 1.505 2.115 1.755 3.245 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 1.115 0.085 1.445 1.13 ;
      RECT 0.115 0.085 0.445 1.01 ;
    LAYER mcon ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_nor2_2

MACRO scs8ls_fah_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 14.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555 1.355 2.895 2.15 ;
        RECT 2.725 0.765 2.895 1.355 ;
        RECT 2.725 0.595 5.435 0.765 ;
        RECT 3.565 0.765 3.735 1.63 ;
        RECT 4.405 0.765 4.595 1.605 ;
        RECT 5.265 0.765 5.435 0.92 ;
        RECT 3.44 1.63 3.77 1.96 ;
        RECT 5.265 0.92 6.205 1.09 ;
        RECT 5.875 1.09 6.205 1.185 ;
    END
    ANTENNAGATEAREA 0.723 ;
  END B

  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.585 1.55 12.92 2.2 ;
        RECT 12.585 0.35 12.835 1.55 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END COUT

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.515 0.8 14.275 1.13 ;
        RECT 13.705 1.13 14.275 1.505 ;
        RECT 13.515 0.355 13.785 0.8 ;
        RECT 13.705 1.505 13.875 1.82 ;
        RECT 13.57 1.82 13.875 2.98 ;
    END
    ANTENNADIFFAREA 0.5618 ;
  END SUM

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.45 1.45 11.875 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END CI

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.29 2.045 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 12.155 0.84 12.325 1.01 ;
      RECT 0.155 1.21 0.325 1.38 ;
      RECT 8.315 0.84 8.485 1.01 ;
      RECT 3.995 1.21 4.165 1.38 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
    LAYER met1 ;
      RECT 8.255 0.995 8.545 1.04 ;
      RECT 8.255 0.855 12.385 0.995 ;
      RECT 12.095 0.995 12.385 1.04 ;
      RECT 8.255 0.81 8.545 0.855 ;
      RECT 12.095 0.81 12.385 0.855 ;
      RECT 0.095 1.365 0.385 1.41 ;
      RECT 0.095 1.225 4.225 1.365 ;
      RECT 3.935 1.365 4.225 1.41 ;
      RECT 0.095 1.18 0.385 1.225 ;
      RECT 3.935 1.18 4.225 1.225 ;
    LAYER li1 ;
      RECT 7.215 2.905 9.575 3.075 ;
      RECT 7.215 2.41 7.385 2.905 ;
      RECT 9.405 1.96 9.575 2.905 ;
      RECT 8.48 1.225 8.735 2.905 ;
      RECT 6.225 2.27 7.385 2.41 ;
      RECT 9.245 1.63 9.575 1.96 ;
      RECT 5.385 2.24 7.385 2.27 ;
      RECT 9.245 0.765 9.415 1.63 ;
      RECT 5.385 2.1 6.395 2.24 ;
      RECT 7.215 1.96 7.385 2.24 ;
      RECT 9.245 0.595 10.255 0.765 ;
      RECT 7.215 1.63 7.505 1.96 ;
      RECT 10.085 0.765 10.255 1.355 ;
      RECT 10.085 1.355 10.47 1.685 ;
      RECT 3.065 1.185 3.235 2.39 ;
      RECT 3.065 0.935 3.395 1.185 ;
      RECT 2.555 2.39 3.45 2.55 ;
      RECT 5.385 2.27 5.555 2.55 ;
      RECT 2.555 2.55 5.555 2.72 ;
      RECT 7.555 2.13 8.31 2.735 ;
      RECT 8.14 1.04 8.31 2.13 ;
      RECT 8.14 0.64 8.555 1.04 ;
      RECT 8.015 0.39 8.555 0.64 ;
      RECT 10.765 0.675 11.865 0.845 ;
      RECT 10.98 0.845 11.865 1.055 ;
      RECT 11.535 0.375 11.865 0.675 ;
      RECT 10.98 1.95 11.93 2.2 ;
      RECT 8.905 2.13 9.235 2.735 ;
      RECT 8.905 1.055 9.075 2.13 ;
      RECT 8.745 0.425 9.075 1.055 ;
      RECT 8.745 0.255 10.935 0.425 ;
      RECT 10.765 0.425 10.935 0.675 ;
      RECT 10.98 1.055 11.24 1.95 ;
      RECT 0.555 1.99 0.885 2.98 ;
      RECT 0.335 1.82 0.885 1.99 ;
      RECT 0.335 1.47 0.65 1.82 ;
      RECT 0.125 1.18 0.65 1.47 ;
      RECT 0.48 1.13 0.65 1.18 ;
      RECT 0.48 0.96 0.965 1.13 ;
      RECT 0.705 0.35 0.965 0.96 ;
      RECT 3.62 2.13 4.11 2.38 ;
      RECT 3.94 1.41 4.11 2.13 ;
      RECT 3.94 1.185 4.235 1.41 ;
      RECT 3.905 0.935 4.235 1.185 ;
      RECT 4.765 1.355 6.545 1.43 ;
      RECT 5.535 1.43 6.545 1.525 ;
      RECT 6.375 1.02 6.545 1.355 ;
      RECT 6.375 0.85 7.005 1.02 ;
      RECT 6.835 0.425 7.005 0.85 ;
      RECT 6.835 0.255 7.845 0.425 ;
      RECT 7.675 0.425 7.845 1.275 ;
      RECT 7.675 1.275 7.97 1.945 ;
      RECT 4.28 2.1 5.215 2.35 ;
      RECT 4.765 1.43 4.935 2.1 ;
      RECT 4.765 0.935 5.095 1.26 ;
      RECT 4.765 1.26 5.705 1.355 ;
      RECT 0 -0.085 14.4 0.085 ;
      RECT 13.955 0.085 14.285 0.63 ;
      RECT 13.015 0.085 13.345 1.13 ;
      RECT 6.335 0.085 6.665 0.68 ;
      RECT 11.105 0.085 11.355 0.505 ;
      RECT 12.075 0.085 12.405 0.64 ;
      RECT 0.17 0.085 0.535 0.79 ;
      RECT 1.875 0.085 2.125 0.845 ;
      RECT 0 3.245 14.4 3.415 ;
      RECT 14.045 1.82 14.295 3.245 ;
      RECT 13.04 2.71 13.37 3.245 ;
      RECT 11.015 2.94 11.395 3.245 ;
      RECT 12.14 2.71 12.47 3.245 ;
      RECT 6.265 2.58 6.595 3.245 ;
      RECT 0.105 2.16 0.36 3.245 ;
      RECT 1.54 1.95 1.87 3.245 ;
      RECT 12.085 0.81 12.415 1.55 ;
      RECT 1.225 0.505 1.705 1.12 ;
      RECT 1.09 1.63 1.34 2.98 ;
      RECT 0.82 1.3 1.395 1.63 ;
      RECT 1.225 1.12 1.395 1.3 ;
      RECT 6.715 1.93 7.045 2.07 ;
      RECT 5.105 1.76 7.045 1.93 ;
      RECT 6.715 1.36 7.045 1.76 ;
      RECT 6.715 1.19 7.505 1.36 ;
      RECT 7.175 0.63 7.505 1.19 ;
      RECT 5.105 1.6 5.365 1.76 ;
      RECT 2.055 2.89 6.055 3.06 ;
      RECT 5.725 2.44 6.055 2.89 ;
      RECT 2.305 0.255 5.935 0.425 ;
      RECT 5.605 0.425 5.935 0.75 ;
      RECT 2.055 2.015 2.385 2.89 ;
      RECT 2.215 1.185 2.385 2.015 ;
      RECT 2.215 1.015 2.555 1.185 ;
      RECT 2.305 0.425 2.555 1.015 ;
      RECT 10.31 2.13 10.81 2.43 ;
      RECT 10.64 1.185 10.81 2.13 ;
      RECT 10.425 1.015 10.81 1.185 ;
      RECT 10.425 0.595 10.595 1.015 ;
      RECT 13.23 1.3 13.535 1.63 ;
      RECT 11.8 2.37 13.4 2.54 ;
      RECT 13.23 1.63 13.4 2.37 ;
      RECT 9.745 2.6 11.97 2.77 ;
      RECT 11.8 2.54 11.97 2.6 ;
      RECT 9.745 2.77 10.075 2.98 ;
      RECT 9.745 2.1 10.075 2.6 ;
      RECT 9.745 1.185 9.915 2.1 ;
      RECT 9.585 0.935 9.915 1.185 ;
  END
END scs8ls_fah_2

MACRO scs8ls_fah_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 15.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.635 1.35 12.98 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END CI

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.51 1.095 1.8 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.675 2.29 5.155 2.91 ;
        RECT 4.675 1.22 4.925 2.29 ;
    END
    ANTENNAGATEAREA 0.723 ;
  END B

  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.96 1.26 11.395 1.85 ;
        RECT 9.89 1.85 11.395 2.1 ;
        RECT 10.96 1.18 11.785 1.26 ;
        RECT 10.475 1.01 11.785 1.18 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END COUT

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.42 2.02 14.755 2.98 ;
        RECT 13.42 1.85 14.755 2.02 ;
        RECT 13.42 2.02 13.75 2.98 ;
        RECT 14.495 1.18 14.745 1.85 ;
        RECT 13.555 1.01 14.745 1.18 ;
        RECT 13.555 0.48 13.805 1.01 ;
        RECT 14.495 0.48 14.745 1.01 ;
    END
    ANTENNADIFFAREA 1.0976 ;
  END SUM

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 15.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 15.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.915 1.58 6.085 1.75 ;
      RECT 9.275 1.58 9.445 1.75 ;
      RECT 3.515 1.95 3.685 2.12 ;
      RECT 3.035 1.58 3.205 1.75 ;
      RECT 3.995 1.58 4.165 1.75 ;
      RECT 5.435 1.58 5.605 1.75 ;
      RECT 6.875 1.95 7.045 2.12 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
    LAYER met1 ;
      RECT 2.975 1.735 3.265 1.78 ;
      RECT 2.975 1.595 5.665 1.735 ;
      RECT 3.935 1.735 4.225 1.78 ;
      RECT 5.375 1.735 5.665 1.78 ;
      RECT 2.975 1.55 3.265 1.595 ;
      RECT 3.935 1.55 4.225 1.595 ;
      RECT 5.375 1.55 5.665 1.595 ;
      RECT 5.855 1.735 6.145 1.78 ;
      RECT 5.855 1.595 9.505 1.735 ;
      RECT 9.215 1.735 9.505 1.78 ;
      RECT 5.855 1.55 6.145 1.595 ;
      RECT 9.215 1.55 9.505 1.595 ;
      RECT 3.455 2.105 3.745 2.15 ;
      RECT 3.455 1.965 7.105 2.105 ;
      RECT 6.815 2.105 7.105 2.15 ;
      RECT 3.455 1.92 3.745 1.965 ;
      RECT 6.815 1.92 7.105 1.965 ;
    LAYER li1 ;
      RECT 3.715 1.55 4.165 1.765 ;
      RECT 3.715 0.63 3.885 1.55 ;
      RECT 5.435 1.375 5.635 1.78 ;
      RECT 5.435 1.09 5.805 1.375 ;
      RECT 6.655 1.405 7.075 2.15 ;
      RECT 8.58 1.9 9.215 2.1 ;
      RECT 9.045 1.775 9.215 1.9 ;
      RECT 9.045 1.55 9.475 1.775 ;
      RECT 9.045 0.935 9.215 1.55 ;
      RECT 5.885 1.55 6.145 1.78 ;
      RECT 5.975 0.875 6.145 1.55 ;
      RECT 5.875 0.595 6.205 0.875 ;
      RECT 0.085 1.17 1.665 1.34 ;
      RECT 1.335 1.34 1.665 1.65 ;
      RECT 0.085 1.97 0.365 2.98 ;
      RECT 0.085 1.34 0.255 1.97 ;
      RECT 0.085 0.35 0.365 1.17 ;
      RECT 9.78 1.35 10.71 1.68 ;
      RECT 6.535 2.49 6.785 2.735 ;
      RECT 6.535 2.32 7.535 2.49 ;
      RECT 7.365 1.285 7.535 2.32 ;
      RECT 7.365 1.105 7.685 1.285 ;
      RECT 7.365 0.935 8.875 1.105 ;
      RECT 8.705 0.765 8.875 0.935 ;
      RECT 8.705 0.595 9.555 0.765 ;
      RECT 9.385 0.765 9.555 1.01 ;
      RECT 9.385 1.01 9.95 1.18 ;
      RECT 9.78 1.18 9.95 1.35 ;
      RECT 8.545 2.61 12.715 2.78 ;
      RECT 12.295 2.78 12.715 2.86 ;
      RECT 12.295 1.95 12.715 2.61 ;
      RECT 12.295 1.01 12.855 1.18 ;
      RECT 12.295 1.18 12.465 1.95 ;
      RECT 6.195 2.905 8.715 3.075 ;
      RECT 8.545 2.78 8.715 2.905 ;
      RECT 6.99 2.725 7.875 2.905 ;
      RECT 6.195 2.15 6.365 2.905 ;
      RECT 7.705 1.65 7.875 2.725 ;
      RECT 6.195 1.98 6.485 2.15 ;
      RECT 7.705 1.48 8.875 1.65 ;
      RECT 6.315 1.215 6.485 1.98 ;
      RECT 8.205 1.32 8.875 1.48 ;
      RECT 6.315 1.045 7.195 1.215 ;
      RECT 6.865 1.015 7.195 1.045 ;
      RECT 4.23 2.46 4.505 2.67 ;
      RECT 2.175 2.29 4.505 2.46 ;
      RECT 4.23 1.935 4.505 2.29 ;
      RECT 2.175 1.79 2.505 2.29 ;
      RECT 4.335 1.31 4.505 1.935 ;
      RECT 2.305 0.625 2.475 1.79 ;
      RECT 4.065 1.045 4.505 1.31 ;
      RECT 1.015 2.8 1.345 2.98 ;
      RECT 1.015 2.63 3.495 2.8 ;
      RECT 3.165 2.8 3.495 2.96 ;
      RECT 1.015 1.97 1.345 2.63 ;
      RECT 1.835 1 2.005 2.63 ;
      RECT 0.975 0.96 2.005 1 ;
      RECT 0.975 0.79 2.135 0.96 ;
      RECT 1.965 0.425 2.135 0.79 ;
      RECT 0.975 0.35 1.305 0.79 ;
      RECT 1.965 0.255 3.415 0.425 ;
      RECT 3.155 0.425 3.415 1.04 ;
      RECT 2.705 1.78 2.96 2.12 ;
      RECT 2.705 1.55 3.205 1.78 ;
      RECT 3.375 1.935 4.03 2.12 ;
      RECT 3.375 1.38 3.545 1.935 ;
      RECT 2.655 1.21 3.545 1.38 ;
      RECT 2.655 0.625 2.985 1.21 ;
      RECT 13.215 1.35 14.325 1.68 ;
      RECT 9.725 0.67 13.385 0.84 ;
      RECT 13.215 0.84 13.385 1.35 ;
      RECT 8.045 2.27 12.125 2.44 ;
      RECT 11.955 0.84 12.125 2.27 ;
      RECT 8.045 2.44 8.375 2.735 ;
      RECT 8.045 2.095 8.375 2.27 ;
      RECT 8.365 0.425 8.535 0.595 ;
      RECT 6.375 0.595 8.535 0.765 ;
      RECT 6.375 0.765 6.705 0.845 ;
      RECT 9.725 0.425 9.895 0.67 ;
      RECT 8.365 0.255 9.895 0.425 ;
      RECT 5.855 2.12 6.025 2.98 ;
      RECT 5.095 1.95 6.025 2.12 ;
      RECT 5.095 0.92 5.265 1.95 ;
      RECT 5.095 0.875 5.405 0.92 ;
      RECT 4.055 0.705 5.405 0.875 ;
      RECT 5.095 0.425 5.405 0.705 ;
      RECT 5.095 0.255 8.195 0.425 ;
      RECT 4.055 0.255 4.385 0.705 ;
      RECT 0 -0.085 15.36 0.085 ;
      RECT 14.915 0.085 15.245 1.26 ;
      RECT 10.965 0.085 11.295 0.5 ;
      RECT 11.965 0.085 12.295 0.5 ;
      RECT 13.035 0.085 13.375 0.5 ;
      RECT 4.585 0.085 4.915 0.535 ;
      RECT 10.065 0.085 10.315 0.5 ;
      RECT 0.545 0.085 0.795 1 ;
      RECT 1.535 0.085 1.795 0.62 ;
      RECT 13.985 0.085 14.315 0.84 ;
      RECT 0 3.245 15.36 3.415 ;
      RECT 14.95 1.82 15.2 3.245 ;
      RECT 11.495 2.95 12.125 3.245 ;
      RECT 12.92 1.95 13.25 3.245 ;
      RECT 9.115 2.95 9.685 3.245 ;
      RECT 5.325 2.29 5.655 3.245 ;
      RECT 1.575 2.97 1.915 3.245 ;
      RECT 0.565 1.97 0.815 3.245 ;
      RECT 10.425 2.95 10.755 3.245 ;
      RECT 13.92 2.19 14.25 3.245 ;
  END
END scs8ls_fah_4

MACRO scs8ls_fahcin_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.515 0.44 12.845 0.84 ;
        RECT 12.595 0.84 12.845 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END SUM

  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.705 1.155 9.035 1.485 ;
    END
    ANTENNAGATEAREA 0.525 ;
  END CIN

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.35 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.875 1.18 5.205 1.585 ;
    END
    ANTENNAGATEAREA 0.723 ;
  END B

  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.64 0.44 8.035 0.985 ;
        RECT 6.64 0.985 7.07 1.31 ;
        RECT 6.9 1.31 7.07 2.335 ;
        RECT 6.82 2.335 7.615 2.665 ;
    END
    ANTENNADIFFAREA 1.9598 ;
  END COUT

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12.96 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12.96 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 4.475 1.95 4.645 2.12 ;
      RECT 2.075 1.95 2.245 2.12 ;
      RECT 7.355 1.95 7.525 2.12 ;
      RECT 10.715 1.95 10.885 2.12 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
    LAYER met1 ;
      RECT 2.015 2.105 2.305 2.15 ;
      RECT 2.015 1.965 10.945 2.105 ;
      RECT 4.415 2.105 4.705 2.15 ;
      RECT 7.295 2.105 7.585 2.15 ;
      RECT 10.655 2.105 10.945 2.15 ;
      RECT 2.015 1.92 2.305 1.965 ;
      RECT 4.415 1.92 4.705 1.965 ;
      RECT 7.295 1.92 7.585 1.965 ;
      RECT 10.655 1.92 10.945 1.965 ;
    LAYER li1 ;
      RECT 1.005 2.905 3.935 3.075 ;
      RECT 3.685 2.25 3.935 2.905 ;
      RECT 1.005 1.63 1.175 2.905 ;
      RECT 1.005 1.3 1.445 1.63 ;
      RECT 1.005 1.18 1.29 1.3 ;
      RECT 0.12 1.01 1.29 1.18 ;
      RECT 1.12 0.425 1.29 1.01 ;
      RECT 1.12 0.255 2.835 0.425 ;
      RECT 2.585 0.425 2.835 0.75 ;
      RECT 0.12 1.18 0.375 2.98 ;
      RECT 0.12 0.35 0.45 1.01 ;
      RECT 9.895 2.57 10.065 2.735 ;
      RECT 9.895 2.4 11.635 2.57 ;
      RECT 11.385 2.57 11.635 2.735 ;
      RECT 9.895 1.9 10.065 2.4 ;
      RECT 11.195 1.85 11.635 2.4 ;
      RECT 11.195 1.25 11.365 1.85 ;
      RECT 11.085 1.22 11.365 1.25 ;
      RECT 11.085 0.66 11.415 1.22 ;
      RECT 0 3.245 12.96 3.415 ;
      RECT 8.885 1.995 9.055 3.245 ;
      RECT 12.145 1.85 12.395 3.245 ;
      RECT 5.405 2.73 5.765 3.245 ;
      RECT 0.575 1.95 0.825 3.245 ;
      RECT 0 -0.085 12.96 0.085 ;
      RECT 8.705 0.085 9.045 0.985 ;
      RECT 11.925 0.085 12.345 0.81 ;
      RECT 0.62 0.085 0.95 0.84 ;
      RECT 5.465 0.085 5.97 0.635 ;
      RECT 1.345 2.565 2.98 2.735 ;
      RECT 2.655 2.045 2.98 2.565 ;
      RECT 1.345 1.82 1.835 2.565 ;
      RECT 2.81 1.09 2.98 2.045 ;
      RECT 1.615 1.02 1.835 1.82 ;
      RECT 2.81 0.92 3.175 1.09 ;
      RECT 1.475 0.615 1.835 1.02 ;
      RECT 3.005 0.425 3.175 0.92 ;
      RECT 3.005 0.255 3.945 0.425 ;
      RECT 3.695 0.425 3.945 1.125 ;
      RECT 2.045 2.07 2.485 2.395 ;
      RECT 2.045 1.89 2.415 2.07 ;
      RECT 2.165 0.615 2.415 1.89 ;
      RECT 7.24 1.17 7.555 2.15 ;
      RECT 10.265 1.26 10.515 2.23 ;
      RECT 10.07 0.74 10.915 1.26 ;
      RECT 10.745 0.49 10.915 0.74 ;
      RECT 10.745 0.32 11.755 0.49 ;
      RECT 11.585 0.49 11.755 1.01 ;
      RECT 11.585 1.01 12.425 1.18 ;
      RECT 12.145 1.18 12.425 1.68 ;
      RECT 4.445 1.875 4.705 2.735 ;
      RECT 4.455 0.67 4.705 1.875 ;
      RECT 5.97 1.82 6.31 2.22 ;
      RECT 6.14 1.065 6.31 1.82 ;
      RECT 6.14 0.385 6.47 1.065 ;
      RECT 8.125 1.82 8.375 2.735 ;
      RECT 8.205 1.065 8.375 1.82 ;
      RECT 8.205 0.385 8.535 1.065 ;
      RECT 9.255 2.905 11.975 3.075 ;
      RECT 10.8 2.74 11.155 2.905 ;
      RECT 9.255 1.995 9.725 2.905 ;
      RECT 11.805 1.68 11.975 2.905 ;
      RECT 9.555 1.34 9.725 1.995 ;
      RECT 11.535 1.35 11.975 1.68 ;
      RECT 9.555 0.74 9.885 1.34 ;
      RECT 10.685 1.43 11.015 2.15 ;
      RECT 4.955 1.99 5.285 2.22 ;
      RECT 4.955 1.82 5.8 1.99 ;
      RECT 5.63 1.585 5.8 1.82 ;
      RECT 5.63 1.255 5.97 1.585 ;
      RECT 5.63 1.01 5.8 1.255 ;
      RECT 4.965 0.84 5.8 1.01 ;
      RECT 4.965 0.425 5.295 0.84 ;
      RECT 4.115 0.255 5.295 0.425 ;
      RECT 4.115 0.425 4.285 1.38 ;
      RECT 3.685 1.38 4.285 1.55 ;
      RECT 3.685 1.55 3.99 1.71 ;
      RECT 6.15 2.905 8.715 3.075 ;
      RECT 8.545 1.825 8.715 2.905 ;
      RECT 8.545 1.655 9.385 1.825 ;
      RECT 9.215 0.57 9.385 1.655 ;
      RECT 9.215 0.255 10.575 0.57 ;
      RECT 7.785 1.485 7.955 2.905 ;
      RECT 7.745 1.155 8.035 1.485 ;
      RECT 4.105 2.905 5.045 3.075 ;
      RECT 4.875 2.56 5.045 2.905 ;
      RECT 4.105 2.05 4.275 2.905 ;
      RECT 3.185 1.88 4.275 2.05 ;
      RECT 3.185 2.05 3.515 2.735 ;
      RECT 3.185 1.875 3.515 1.88 ;
      RECT 3.345 0.595 3.515 1.875 ;
      RECT 4.875 2.39 6.65 2.56 ;
      RECT 6.15 2.56 6.65 2.905 ;
      RECT 6.48 1.84 6.65 2.39 ;
      RECT 6.48 1.51 6.73 1.84 ;
  END
END scs8ls_fahcin_1

MACRO scs8ls_fahcon_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 11.52 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN COUTN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.32 0.35 6.65 1.21 ;
        RECT 6.005 1.21 6.65 1.38 ;
        RECT 6.005 1.38 6.175 2.085 ;
        RECT 5.79 2.085 6.175 2.255 ;
        RECT 5.79 2.255 6.12 2.965 ;
    END
    ANTENNADIFFAREA 0.7826 ;
  END COUTN

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.075 1.82 11.435 2.98 ;
        RECT 11.265 1.13 11.435 1.82 ;
        RECT 11.155 0.35 11.435 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END SUM

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.35 0.805 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.18 5.06 1.55 ;
    END
    ANTENNAGATEAREA 0.969 ;
  END B

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.675 1.18 8.005 1.55 ;
    END
    ANTENNAGATEAREA 0.525 ;
  END CI

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.52 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.52 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 9.275 0.84 9.445 1.01 ;
      RECT 6.875 0.84 7.045 1.01 ;
      RECT 8.795 1.58 8.965 1.75 ;
      RECT 3.035 1.58 3.205 1.75 ;
      RECT 5.915 0.84 6.085 1.01 ;
      RECT 6.395 1.58 6.565 1.75 ;
      RECT 2.075 0.84 2.245 1.01 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
    LAYER met1 ;
      RECT 2.975 1.735 3.265 1.78 ;
      RECT 2.975 1.595 9.025 1.735 ;
      RECT 6.335 1.735 6.625 1.78 ;
      RECT 8.735 1.735 9.025 1.78 ;
      RECT 2.975 1.55 3.265 1.595 ;
      RECT 6.335 1.55 6.625 1.595 ;
      RECT 8.735 1.55 9.025 1.595 ;
      RECT 2.015 0.995 2.305 1.04 ;
      RECT 2.015 0.855 9.505 0.995 ;
      RECT 5.855 0.995 6.145 1.04 ;
      RECT 6.815 0.995 7.105 1.04 ;
      RECT 9.215 0.995 9.505 1.04 ;
      RECT 2.015 0.81 2.305 0.855 ;
      RECT 5.855 0.81 6.145 0.855 ;
      RECT 6.815 0.81 7.105 0.855 ;
      RECT 9.215 0.81 9.505 0.855 ;
    LAYER li1 ;
      RECT 0 3.245 11.52 3.415 ;
      RECT 10.65 2.1 10.9 3.245 ;
      RECT 7.645 1.94 7.815 3.245 ;
      RECT 0.655 1.95 0.985 3.245 ;
      RECT 4.545 1.805 4.875 3.245 ;
      RECT 0 -0.085 11.52 0.085 ;
      RECT 7.745 0.085 7.995 1.01 ;
      RECT 10.495 0.085 10.895 0.41 ;
      RECT 0.545 0.48 0.905 0.81 ;
      RECT 0.545 0.085 0.715 0.48 ;
      RECT 4.905 0.085 5.155 0.965 ;
      RECT 8.515 1.55 8.965 1.78 ;
      RECT 8.515 1.3 8.765 1.55 ;
      RECT 6.345 1.55 6.61 1.88 ;
      RECT 6.345 2.085 7.475 2.97 ;
      RECT 7.305 0.96 7.475 2.085 ;
      RECT 7.245 0.35 7.575 0.96 ;
      RECT 6.82 1.13 7.135 1.8 ;
      RECT 6.82 0.81 7.075 1.13 ;
      RECT 8.575 2.87 10.455 3.04 ;
      RECT 8.575 2.66 8.905 2.87 ;
      RECT 10.2 1.93 10.455 2.87 ;
      RECT 10.2 1.76 10.625 1.93 ;
      RECT 10.455 1.09 10.625 1.76 ;
      RECT 9.815 0.92 10.625 1.09 ;
      RECT 9.815 0.595 9.985 0.92 ;
      RECT 4.04 0.425 4.735 1.01 ;
      RECT 2.785 0.255 4.735 0.425 ;
      RECT 4.04 1.805 4.375 2.965 ;
      RECT 4.04 1.01 4.21 1.805 ;
      RECT 2.785 0.425 3.115 0.555 ;
      RECT 9.475 1.26 9.69 1.59 ;
      RECT 9.475 1.04 9.645 1.26 ;
      RECT 9.275 0.81 9.645 1.04 ;
      RECT 5.665 0.81 6.115 1.04 ;
      RECT 5.57 1.475 5.835 1.805 ;
      RECT 5.665 1.04 5.835 1.475 ;
      RECT 10.81 1.3 11.095 1.63 ;
      RECT 9.135 1.82 9.36 2.15 ;
      RECT 9.135 1.38 9.305 1.82 ;
      RECT 8.935 1.21 9.305 1.38 ;
      RECT 8.935 1.13 9.105 1.21 ;
      RECT 8.775 0.425 9.105 1.13 ;
      RECT 8.775 0.255 10.325 0.425 ;
      RECT 10.155 0.425 10.325 0.58 ;
      RECT 10.155 0.58 10.98 0.75 ;
      RECT 10.81 0.75 10.98 1.3 ;
      RECT 2.03 2.225 3.275 2.395 ;
      RECT 2.03 2 2.2 2.225 ;
      RECT 2.945 0.725 3.275 2.225 ;
      RECT 0.085 1.95 0.485 2.98 ;
      RECT 0.085 1.15 1.18 1.18 ;
      RECT 0.975 1.18 1.18 1.68 ;
      RECT 0.085 0.98 1.245 1.15 ;
      RECT 1.075 0.425 1.245 0.98 ;
      RECT 1.075 0.255 2.615 0.425 ;
      RECT 2.445 0.425 2.615 0.725 ;
      RECT 2.445 0.725 2.775 1.805 ;
      RECT 2.4 1.805 2.775 2.055 ;
      RECT 0.085 1.18 0.255 1.95 ;
      RECT 0.085 0.48 0.365 0.98 ;
      RECT 1.19 2.905 3.81 3.075 ;
      RECT 1.19 1.85 1.52 2.905 ;
      RECT 3.46 0.645 3.81 2.905 ;
      RECT 1.35 1.49 1.52 1.85 ;
      RECT 1.35 1.32 1.745 1.49 ;
      RECT 1.415 0.595 1.745 1.32 ;
      RECT 5.325 0.39 6.15 0.64 ;
      RECT 5.1 1.975 5.43 2.965 ;
      RECT 5.23 1.305 5.4 1.975 ;
      RECT 5.23 1.135 5.495 1.305 ;
      RECT 5.325 0.64 5.495 1.135 ;
      RECT 8.015 2.49 8.345 2.98 ;
      RECT 8.015 2.32 10.03 2.49 ;
      RECT 9.56 2.49 10.03 2.7 ;
      RECT 8.015 1.82 8.345 2.32 ;
      RECT 9.56 1.82 10.03 2.32 ;
      RECT 8.175 1.13 8.345 1.82 ;
      RECT 9.86 1.59 10.03 1.82 ;
      RECT 8.175 0.35 8.515 1.13 ;
      RECT 9.86 1.26 10.285 1.59 ;
      RECT 1.69 2.565 3.26 2.735 ;
      RECT 1.69 1.83 1.86 2.565 ;
      RECT 1.69 1.66 2.095 1.83 ;
      RECT 1.925 1.325 2.095 1.66 ;
      RECT 1.925 0.595 2.275 1.325 ;
  END
END scs8ls_fahcon_1

MACRO scs8ls_fill_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.48 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.48 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.48 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 0.48 0.085 ;
      RECT 0 3.245 0.48 3.415 ;
    LAYER mcon ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_fill_1

MACRO scs8ls_fill_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.96 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.96 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 0.96 0.085 ;
      RECT 0 3.245 0.96 3.415 ;
    LAYER mcon ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_fill_2

MACRO scs8ls_fill_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.92 0.085 ;
      RECT 0 3.245 1.92 3.415 ;
    LAYER mcon ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
  END
END scs8ls_fill_4

MACRO scs8ls_fill_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 0 3.245 3.84 3.415 ;
    LAYER mcon ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
  END
END scs8ls_fill_8

MACRO scs8ls_ha_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.45 0.255 2.78 0.67 ;
    END
    ANTENNAGATEAREA 0.468 ;
  END A

  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.31 1.85 4.715 2.98 ;
        RECT 4.545 1.18 4.715 1.85 ;
        RECT 4.31 0.475 4.715 1.18 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END COUT

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.35 0.445 1.13 ;
        RECT 0.115 1.13 0.355 1.82 ;
        RECT 0.115 1.82 0.445 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END SUM

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.765 1.55 3.3 1.8 ;
        RECT 1.765 1.47 2.095 1.55 ;
        RECT 2.97 1.47 3.3 1.55 ;
    END
    ANTENNAGATEAREA 0.468 ;
  END B

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.47 1.35 4.375 1.68 ;
      RECT 3.36 2.14 3.64 2.98 ;
      RECT 1.195 1.97 3.64 2.14 ;
      RECT 3.47 1.68 3.64 1.97 ;
      RECT 3.47 1.255 3.64 1.35 ;
      RECT 3.02 1.085 3.64 1.255 ;
      RECT 3.02 0.575 3.35 1.085 ;
      RECT 1.195 1.47 1.525 1.97 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 3.81 0.085 4.14 1.18 ;
      RECT 0.625 0.085 0.875 0.795 ;
      RECT 1.93 0.085 2.28 0.96 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 0.615 2.65 1.205 3.245 ;
      RECT 2.485 2.31 3.19 3.245 ;
      RECT 3.81 2.1 4.14 3.245 ;
      RECT 1.41 2.48 1.74 2.8 ;
      RECT 0.685 2.31 1.74 2.48 ;
      RECT 0.685 1.63 0.855 2.31 ;
      RECT 0.525 1.3 0.855 1.63 ;
      RECT 0.685 1.13 1.4 1.3 ;
      RECT 1.07 0.91 1.4 1.13 ;
      RECT 2.46 1.3 2.79 1.355 ;
      RECT 1.58 1.13 2.79 1.3 ;
      RECT 2.46 0.84 2.79 1.13 ;
      RECT 1.58 0.63 1.75 1.13 ;
    LAYER mcon ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_ha_1

MACRO scs8ls_ha_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.885 0.35 5.215 1.13 ;
        RECT 4.885 1.13 5.055 1.82 ;
        RECT 4.865 1.82 5.195 2.17 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END COUT

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.82 4.675 2.17 ;
        RECT 4.505 1.05 4.675 1.82 ;
        RECT 3.975 0.88 4.675 1.05 ;
    END
    ANTENNADIFFAREA 0.5802 ;
  END SUM

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.06 1.45 1.39 1.78 ;
    END
    ANTENNAGATEAREA 0.522 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 2.32 2.12 2.52 ;
        RECT 0.125 1.63 0.295 2.32 ;
        RECT 1.79 1.45 2.12 2.32 ;
        RECT 0.125 1.3 0.55 1.63 ;
    END
    ANTENNAGATEAREA 0.522 ;
  END B

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 5.395 0.085 5.645 1.13 ;
      RECT 4.455 0.085 4.705 0.71 ;
      RECT 0.935 0.085 1.265 0.6 ;
      RECT 1.795 0.085 2.125 0.6 ;
      RECT 3.545 0.085 3.875 0.71 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 0.115 2.69 0.445 3.245 ;
      RECT 1.015 2.69 1.4 3.245 ;
      RECT 3.08 2.68 3.845 3.245 ;
      RECT 4.415 2.68 4.745 3.245 ;
      RECT 5.315 2.68 5.645 3.245 ;
      RECT 3.32 1.22 4.33 1.55 ;
      RECT 2.63 1.92 3.49 2.17 ;
      RECT 3.32 1.55 3.49 1.92 ;
      RECT 3.32 1.11 3.49 1.22 ;
      RECT 2.635 0.94 3.49 1.11 ;
      RECT 2.635 0.595 2.805 0.94 ;
      RECT 1.365 0.77 2.465 0.94 ;
      RECT 2.295 0.425 2.465 0.77 ;
      RECT 2.295 0.255 3.315 0.425 ;
      RECT 2.985 0.425 3.315 0.77 ;
      RECT 2.29 2.34 5.555 2.51 ;
      RECT 5.385 1.63 5.555 2.34 ;
      RECT 5.225 1.3 5.555 1.63 ;
      RECT 2.29 1.61 2.46 2.34 ;
      RECT 2.29 1.28 3.035 1.61 ;
      RECT 0.72 1.13 2.46 1.28 ;
      RECT 0.115 1.11 2.46 1.13 ;
      RECT 0.72 1.28 0.89 1.98 ;
      RECT 0.565 1.98 0.895 2.15 ;
      RECT 0.115 0.96 0.89 1.11 ;
      RECT 0.115 0.35 0.445 0.96 ;
    LAYER mcon ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_ha_2

MACRO scs8ls_ha_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.455 1.315 1.785 ;
    END
    ANTENNAGATEAREA 0.936 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.455 2.275 1.785 ;
    END
    ANTENNAGATEAREA 0.936 ;
  END B

  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.21 1.13 7.555 1.82 ;
        RECT 6.22 1.82 7.555 2.15 ;
        RECT 6.35 0.88 7.555 1.13 ;
        RECT 6.35 0.35 6.6 0.88 ;
    END
    ANTENNADIFFAREA 1.2656 ;
  END COUT

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
    END
  END vpwr

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 8.735 1.965 9.985 2.105 ;
        RECT 9.695 2.105 9.985 2.15 ;
        RECT 9.695 1.92 9.985 1.965 ;
        RECT 8.735 2.105 9.025 2.15 ;
        RECT 8.735 1.92 9.025 1.965 ;
    END
    ANTENNADIFFAREA 1.4701 ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met1 ;
  END SUM

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 10.08 0.085 ;
      RECT 7.64 0.085 7.97 0.71 ;
      RECT 8.57 0.085 8.9 0.81 ;
      RECT 9.58 0.085 9.885 0.81 ;
      RECT 0.545 0.085 0.795 0.945 ;
      RECT 1.41 0.085 1.66 0.945 ;
      RECT 4.95 0.085 5.28 1.255 ;
      RECT 5.92 0.085 6.17 1.13 ;
      RECT 6.78 0.085 7.11 0.71 ;
      RECT 3.9 2.335 7.895 2.49 ;
      RECT 3.085 2.32 7.895 2.335 ;
      RECT 7.725 1.65 7.895 2.32 ;
      RECT 7.725 1.32 9.645 1.65 ;
      RECT 3.085 2.235 4.07 2.32 ;
      RECT 2.925 2.165 4.07 2.235 ;
      RECT 2.925 2.125 3.255 2.165 ;
      RECT 1.455 1.955 3.255 2.125 ;
      RECT 1.455 2.125 1.735 2.735 ;
      RECT 2.5 1.905 3.255 1.955 ;
      RECT 2.5 1.285 2.67 1.905 ;
      RECT 2.34 0.605 2.67 1.285 ;
      RECT 8.075 2.15 8.305 2.98 ;
      RECT 8.075 1.82 9.995 2.15 ;
      RECT 9.075 2.15 9.405 2.98 ;
      RECT 9.825 1.15 9.995 1.82 ;
      RECT 8.15 0.98 9.995 1.15 ;
      RECT 8.15 0.35 8.4 0.98 ;
      RECT 9.07 0.35 9.4 0.98 ;
      RECT 5.88 1.32 6.955 1.65 ;
      RECT 4.955 1.995 6.05 2.15 ;
      RECT 3.9 1.82 6.05 1.995 ;
      RECT 3.9 1.745 4.23 1.82 ;
      RECT 5.88 1.65 6.05 1.82 ;
      RECT 3.9 1.735 4.07 1.745 ;
      RECT 3.075 1.575 4.07 1.735 ;
      RECT 3.075 1.405 4.28 1.575 ;
      RECT 3.95 0.655 4.28 1.405 ;
      RECT 0 3.245 10.08 3.415 ;
      RECT 4.43 2.66 4.76 3.245 ;
      RECT 5.49 2.66 5.945 3.245 ;
      RECT 6.675 2.66 7.005 3.245 ;
      RECT 7.575 2.66 7.905 3.245 ;
      RECT 3.375 2.505 3.705 3.245 ;
      RECT 2.475 2.405 2.805 3.245 ;
      RECT 8.475 2.32 8.805 3.245 ;
      RECT 9.635 2.32 9.965 3.245 ;
      RECT 0.555 2.295 0.805 3.245 ;
      RECT 4.45 1.425 5.71 1.595 ;
      RECT 5.46 0.575 5.71 1.425 ;
      RECT 4.45 0.485 4.78 1.425 ;
      RECT 3.52 0.315 4.78 0.485 ;
      RECT 3.52 0.485 3.78 1.235 ;
      RECT 0.115 1.115 2.17 1.285 ;
      RECT 0.115 0.605 0.365 1.115 ;
      RECT 0.98 0.605 1.23 1.115 ;
      RECT 1.84 0.435 2.17 1.115 ;
      RECT 1.84 0.265 3.17 0.435 ;
      RECT 2.84 0.435 3.17 1.235 ;
      RECT 1.005 2.905 2.235 3.075 ;
      RECT 1.905 2.295 2.235 2.905 ;
      RECT 1.005 2.125 1.255 2.905 ;
      RECT 0.105 1.955 1.255 2.125 ;
      RECT 0.105 2.125 0.385 2.965 ;
    LAYER mcon ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 1.95 9.925 2.12 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 1.95 8.965 2.12 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_ha_4

MACRO scs8ls_inv_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.3 0.815 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985 0.35 1.315 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 1.44 3.415 ;
      RECT 0.485 1.95 0.815 3.245 ;
      RECT 0 -0.085 1.44 0.085 ;
      RECT 0.485 0.085 0.815 1.13 ;
    LAYER mcon ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_inv_1

MACRO scs8ls_inv_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.085 1.55 7.07 1.78 ;
    END
    ANTENNAGATEAREA 4.464 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.585 1.92 7.575 2.15 ;
    END
    ANTENNADIFFAREA 4.3792 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 1.055 1.94 1.345 3.245 ;
      RECT 2.045 1.94 2.295 3.245 ;
      RECT 2.995 1.94 3.245 3.245 ;
      RECT 3.915 1.94 4.15 3.245 ;
      RECT 4.81 1.94 5.095 3.245 ;
      RECT 5.765 1.94 6.095 3.245 ;
      RECT 6.765 1.94 7.095 3.245 ;
      RECT 0.115 1.82 0.365 3.245 ;
      RECT 7.735 1.82 8.045 3.245 ;
      RECT 7.265 1.13 7.545 2.98 ;
      RECT 7.215 0.35 7.545 1.13 ;
      RECT 6.265 1.285 6.595 2.98 ;
      RECT 6.265 1.18 6.525 1.285 ;
      RECT 6.195 0.35 6.525 1.18 ;
      RECT 5.265 1.285 5.58 2.98 ;
      RECT 5.265 1.18 5.525 1.285 ;
      RECT 5.215 0.35 5.525 1.18 ;
      RECT 4.34 1.94 4.63 2.98 ;
      RECT 4.34 0.35 4.595 1.94 ;
      RECT 3.415 0.35 3.71 2.98 ;
      RECT 2.465 1.94 2.795 2.98 ;
      RECT 2.485 0.35 2.795 1.94 ;
      RECT 1.07 1.35 1.38 1.77 ;
      RECT 2.02 1.35 2.31 1.77 ;
      RECT 2.97 1.35 3.245 1.77 ;
      RECT 3.885 1.35 4.165 1.77 ;
      RECT 4.77 1.35 5.085 1.77 ;
      RECT 5.755 1.35 6.09 1.77 ;
      RECT 6.77 1.35 7.09 1.77 ;
      RECT 1.515 1.94 1.845 2.98 ;
      RECT 1.555 0.35 1.845 1.94 ;
      RECT 0.565 1.33 0.885 2.995 ;
      RECT 0.615 1.13 0.885 1.33 ;
      RECT 0.615 0.35 0.945 1.13 ;
      RECT 0.185 0.085 0.445 1.13 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 1.115 0.085 1.375 1.13 ;
      RECT 2.025 0.085 2.305 1.13 ;
      RECT 2.975 0.085 3.245 1.13 ;
      RECT 3.89 0.085 4.15 1.13 ;
      RECT 4.765 0.085 5.025 1.13 ;
      RECT 5.705 0.085 6.025 1.13 ;
      RECT 6.705 0.085 7.045 1.13 ;
      RECT 7.715 0.085 8.045 1.13 ;
    LAYER mcon ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 0.645 1.95 0.815 2.12 ;
      RECT 1.595 1.95 1.765 2.12 ;
      RECT 2.545 1.95 2.715 2.12 ;
      RECT 3.495 1.95 3.665 2.12 ;
      RECT 4.395 1.95 4.565 2.12 ;
      RECT 5.345 1.95 5.515 2.12 ;
      RECT 6.345 1.95 6.515 2.12 ;
      RECT 7.345 1.95 7.515 2.12 ;
      RECT 6.84 1.58 7.01 1.75 ;
      RECT 5.845 1.58 6.015 1.75 ;
      RECT 4.85 1.58 5.02 1.75 ;
      RECT 3.94 1.58 4.11 1.75 ;
      RECT 3.025 1.58 3.195 1.75 ;
      RECT 2.085 1.58 2.255 1.75 ;
      RECT 1.145 1.58 1.315 1.75 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
  END
END scs8ls_inv_16

MACRO scs8ls_inv_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.56 0.35 0.89 1.13 ;
        RECT 0.605 1.13 0.89 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.3 0.435 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 1.44 3.415 ;
      RECT 1.085 1.82 1.335 3.245 ;
      RECT 0.105 1.95 0.435 3.245 ;
      RECT 0 -0.085 1.44 0.085 ;
      RECT 1.07 0.085 1.32 1.13 ;
      RECT 0.13 0.085 0.38 1.13 ;
    LAYER mcon ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_inv_2

MACRO scs8ls_inv_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.8 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.18 2.275 1.95 ;
        RECT 0.6 1.95 2.275 2.12 ;
        RECT 0.615 1.01 2.275 1.18 ;
        RECT 0.6 2.12 0.93 2.98 ;
        RECT 1.5 2.12 1.83 2.98 ;
        RECT 0.615 0.35 0.865 1.01 ;
        RECT 1.605 0.35 1.775 1.01 ;
    END
    ANTENNADIFFAREA 1.116 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 2.4 3.415 ;
      RECT 2.03 2.29 2.28 3.245 ;
      RECT 0.15 1.95 0.4 3.245 ;
      RECT 1.13 2.29 1.3 3.245 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 1.955 0.085 2.285 0.84 ;
      RECT 0.115 0.085 0.445 1.13 ;
      RECT 1.045 0.085 1.375 0.84 ;
    LAYER mcon ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_inv_4

MACRO scs8ls_inv_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.42 1.18 4.195 1.31 ;
        RECT 2.495 1.31 4.195 1.62 ;
        RECT 0.56 1.14 4.195 1.18 ;
        RECT 2.495 1.62 2.665 1.95 ;
        RECT 3.365 1.62 3.695 2.98 ;
        RECT 0.56 1.01 2.68 1.14 ;
        RECT 3.35 0.35 3.61 1.14 ;
        RECT 0.565 1.95 2.665 2.12 ;
        RECT 0.56 0.35 0.81 1.01 ;
        RECT 1.5 0.35 1.67 1.01 ;
        RECT 2.35 0.35 2.68 1.01 ;
        RECT 0.565 2.12 0.815 2.98 ;
        RECT 1.515 2.12 1.845 2.98 ;
        RECT 2.495 2.12 2.665 2.98 ;
    END
    ANTENNADIFFAREA 2.1728 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.56 1.35 2.25 1.78 ;
    END
    ANTENNAGATEAREA 2.232 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 3.78 0.085 4.11 0.97 ;
      RECT 0.13 0.085 0.38 1.13 ;
      RECT 0.99 0.085 1.32 0.84 ;
      RECT 1.85 0.085 2.18 0.84 ;
      RECT 2.85 0.085 3.18 0.97 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 3.865 1.82 4.195 3.245 ;
      RECT 0.115 1.82 0.365 3.245 ;
      RECT 1.015 2.29 1.345 3.245 ;
      RECT 2.045 2.29 2.295 3.245 ;
      RECT 2.865 1.82 3.195 3.245 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_inv_8

MACRO scs8ls_maj3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.285 1.43 3.575 1.76 ;
        RECT 2.285 1.76 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END C

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.85 0.49 2.98 ;
        RECT 0.085 1.18 0.255 1.85 ;
        RECT 0.085 0.48 0.445 1.18 ;
    END
    ANTENNADIFFAREA 0.5385 ;
  END X

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.43 1.685 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.645 0.255 3.715 0.57 ;
        RECT 3.485 0.57 3.715 0.67 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.565 1.95 3.725 2.12 ;
      RECT 3.395 2.12 3.725 2.94 ;
      RECT 3.395 1.93 3.725 1.95 ;
      RECT 0.615 1.09 3.7 1.26 ;
      RECT 3.37 0.84 3.7 1.09 ;
      RECT 1.565 2.12 1.895 2.94 ;
      RECT 1.895 1.26 2.065 1.95 ;
      RECT 1.48 0.58 1.81 1.09 ;
      RECT 0.615 1.26 0.785 1.35 ;
      RECT 0.425 1.35 0.785 1.68 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 2.305 0.085 2.475 0.74 ;
      RECT 0.615 0.085 0.99 0.91 ;
      RECT 2.305 0.74 2.85 0.91 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 2.435 2.29 2.84 3.245 ;
      RECT 0.66 1.95 0.99 3.245 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_maj3_1

MACRO scs8ls_maj3_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.18 1.795 1.55 ;
    END
    ANTENNAGATEAREA 0.522 ;
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555 1.82 0.915 2.98 ;
        RECT 0.555 1.13 0.725 1.82 ;
        RECT 0.555 0.35 0.895 1.13 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.215 1.63 3.715 1.78 ;
        RECT 3.215 1.3 4.535 1.63 ;
        RECT 3.215 1.245 3.715 1.3 ;
    END
    ANTENNAGATEAREA 0.522 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.305 1.245 2.975 1.78 ;
    END
    ANTENNAGATEAREA 0.522 ;
  END B

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.965 1.95 4.685 2.12 ;
      RECT 4.355 2.12 4.685 2.86 ;
      RECT 4.355 1.82 4.685 1.95 ;
      RECT 1.965 0.905 4.66 1.075 ;
      RECT 4.33 1.075 4.66 1.13 ;
      RECT 4.33 0.35 4.66 0.905 ;
      RECT 1.965 2.12 2.785 2.755 ;
      RECT 1.965 0.35 2.76 0.905 ;
      RECT 1.085 1.78 2.135 1.95 ;
      RECT 1.965 1.075 2.135 1.78 ;
      RECT 1.085 1.65 1.255 1.78 ;
      RECT 0.895 1.32 1.255 1.65 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 3.485 2.29 3.815 3.245 ;
      RECT 1.085 2.12 1.78 3.245 ;
      RECT 0.135 1.82 0.385 3.245 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 1.075 0.085 1.795 1.01 ;
      RECT 3.34 0.085 3.84 0.68 ;
      RECT 0.135 0.085 0.385 1.13 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_maj3_2

MACRO scs8ls_maj3_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.8 1.47 2.275 1.8 ;
        RECT 2.105 1.8 2.275 1.875 ;
        RECT 2.105 1.875 4.57 2.045 ;
        RECT 4.24 1.47 4.57 1.875 ;
    END
    ANTENNAGATEAREA 0.984 ;
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805 1.175 8.035 1.48 ;
        RECT 7.345 1.48 8.035 1.65 ;
        RECT 6.425 1.005 8.035 1.175 ;
        RECT 7.345 1.65 7.515 1.845 ;
        RECT 6.425 0.475 6.675 1.005 ;
        RECT 6.365 1.845 7.515 2.015 ;
        RECT 6.365 2.015 6.695 2.98 ;
        RECT 7.345 2.015 7.515 2.98 ;
    END
    ANTENNADIFFAREA 1.116 ;
  END X

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.135 1.13 3.235 1.3 ;
        RECT 1.135 1.3 1.465 1.705 ;
        RECT 2.525 1.3 3.235 1.705 ;
    END
    ANTENNAGATEAREA 0.984 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.13 4.925 1.3 ;
        RECT 4.755 1.3 4.925 1.47 ;
        RECT 3.485 1.3 4.01 1.705 ;
        RECT 4.755 1.47 5.22 1.8 ;
    END
    ANTENNAGATEAREA 0.984 ;
  END C

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.58 2.905 1.86 3.075 ;
      RECT 1.53 2.555 1.86 2.905 ;
      RECT 0.58 2.215 0.91 2.905 ;
      RECT 2.49 2.905 3.82 3.075 ;
      RECT 2.49 2.555 2.82 2.905 ;
      RECT 3.49 2.555 3.82 2.905 ;
      RECT 4.51 2.725 4.84 2.98 ;
      RECT 4.51 2.555 5.74 2.725 ;
      RECT 5.41 2.725 5.74 2.98 ;
      RECT 0.625 0.435 0.955 0.62 ;
      RECT 0.625 0.265 1.965 0.435 ;
      RECT 1.635 0.435 1.965 0.96 ;
      RECT 4.505 0.425 4.835 0.62 ;
      RECT 4.505 0.255 5.775 0.425 ;
      RECT 5.445 0.425 5.775 0.96 ;
      RECT 5.39 1.345 7.15 1.675 ;
      RECT 1.095 2.215 5.29 2.385 ;
      RECT 4.96 2.14 5.29 2.215 ;
      RECT 4.96 1.97 5.56 2.14 ;
      RECT 5.39 1.675 5.56 1.97 ;
      RECT 5.39 1.3 5.56 1.345 ;
      RECT 5.095 1.13 5.56 1.3 ;
      RECT 5.095 0.96 5.265 1.13 ;
      RECT 3.065 0.79 5.265 0.96 ;
      RECT 5.095 0.595 5.265 0.79 ;
      RECT 0.795 0.96 0.965 1.875 ;
      RECT 1.095 2.385 1.35 2.735 ;
      RECT 1.095 2.045 1.41 2.215 ;
      RECT 0.795 1.875 1.41 2.045 ;
      RECT 0.795 0.79 1.465 0.96 ;
      RECT 1.135 0.605 1.465 0.79 ;
      RECT 2.99 2.385 3.32 2.735 ;
      RECT 3.065 0.605 3.315 0.79 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 7.715 0.085 8.045 0.835 ;
      RECT 4.005 0.085 4.335 0.62 ;
      RECT 5.955 0.085 6.205 1.175 ;
      RECT 6.855 0.085 7.185 0.835 ;
      RECT 2.145 0.085 2.315 0.96 ;
      RECT 0.115 0.085 0.445 1.285 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 7.715 1.82 8.045 3.245 ;
      RECT 3.99 2.555 4.32 3.245 ;
      RECT 5.94 1.94 6.19 3.245 ;
      RECT 6.895 2.185 7.145 3.245 ;
      RECT 0.13 1.94 0.38 3.245 ;
      RECT 2.06 2.555 2.32 3.245 ;
      RECT 2.495 0.435 2.885 0.935 ;
      RECT 2.495 0.265 3.825 0.435 ;
      RECT 3.495 0.435 3.825 0.62 ;
    LAYER mcon ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
  END
END scs8ls_maj3_4

MACRO scs8ls_mux2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515 0.81 2.785 0.98 ;
        RECT 2.455 0.98 2.785 1.55 ;
        RECT 1.515 0.98 1.685 1.22 ;
        RECT 1.345 1.22 1.685 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885 1.18 2.275 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A0

  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.505 1.35 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.47 ;
  END S

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.795 1.82 4.235 2.98 ;
        RECT 4.065 1.13 4.235 1.82 ;
        RECT 3.865 0.35 4.235 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 3.295 0.085 3.625 0.81 ;
      RECT 0.625 0.68 0.835 1.13 ;
      RECT 0.625 0.085 1.005 0.68 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 0.65 2.4 0.98 3.245 ;
      RECT 3.295 1.82 3.625 3.245 ;
      RECT 3.525 1.3 3.895 1.63 ;
      RECT 1.175 0.39 3.125 0.64 ;
      RECT 2.955 0.64 3.125 0.98 ;
      RECT 2.955 0.98 3.695 1.15 ;
      RECT 3.525 1.15 3.695 1.3 ;
      RECT 2.065 1.89 2.395 2.735 ;
      RECT 1.005 1.72 2.395 1.89 ;
      RECT 1.005 1.02 1.175 1.72 ;
      RECT 1.005 0.85 1.345 1.02 ;
      RECT 1.175 0.64 1.345 0.85 ;
      RECT 1.15 2.905 3.125 3.075 ;
      RECT 2.955 1.65 3.125 2.905 ;
      RECT 2.955 1.32 3.355 1.65 ;
      RECT 1.15 2.23 1.32 2.905 ;
      RECT 0.115 2.06 1.32 2.23 ;
      RECT 0.115 2.23 0.445 2.7 ;
      RECT 0.115 1.95 0.445 2.06 ;
      RECT 0.115 1.13 0.285 1.95 ;
      RECT 0.115 0.54 0.445 1.13 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_mux2_1

MACRO scs8ls_mux2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 0.77 4.665 2.14 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.435 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.18 1.195 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.715 1.45 2.385 1.78 ;
        RECT 2.215 1.3 2.385 1.45 ;
        RECT 2.215 1.13 3.455 1.3 ;
        RECT 3.125 1.3 3.455 1.46 ;
    END
    ANTENNAGATEAREA 0.47 ;
  END S

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 5.28 3.415 ;
      RECT 2.075 2.65 2.405 3.245 ;
      RECT 3.87 2.65 4.21 3.245 ;
      RECT 4.78 2.65 5.165 3.245 ;
      RECT 2.995 2.31 5.165 2.48 ;
      RECT 4.835 1.3 5.165 2.31 ;
      RECT 0.62 1.97 3.165 2.14 ;
      RECT 2.995 2.14 3.165 2.31 ;
      RECT 0.62 2.14 0.84 2.725 ;
      RECT 0.62 1.82 1.535 1.97 ;
      RECT 1.365 1.01 1.535 1.82 ;
      RECT 0.67 0.68 1.535 1.01 ;
      RECT 3.335 1.8 3.795 2.14 ;
      RECT 2.555 1.63 3.795 1.8 ;
      RECT 3.625 0.94 3.795 1.63 ;
      RECT 3.34 0.77 3.795 0.94 ;
      RECT 3.34 0.35 3.67 0.77 ;
      RECT 2.555 1.47 2.885 1.63 ;
      RECT 1.015 2.48 1.345 2.735 ;
      RECT 1.015 2.31 2.825 2.48 ;
      RECT 2.575 2.48 2.825 2.98 ;
      RECT 0.17 0.46 0.5 1.01 ;
      RECT 0.17 0.29 2.75 0.46 ;
      RECT 2.42 0.46 2.75 0.62 ;
      RECT 0 -0.085 5.28 0.085 ;
      RECT 3.84 0.085 4.23 0.6 ;
      RECT 4.835 0.085 5.165 1.13 ;
      RECT 1.715 0.96 2.045 1.13 ;
      RECT 1.715 0.79 3.17 0.96 ;
      RECT 3 0.085 3.17 0.79 ;
      RECT 0.115 2.905 1.905 3.075 ;
      RECT 1.575 2.65 1.905 2.905 ;
      RECT 0.115 1.825 0.445 2.905 ;
    LAYER mcon ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
  END
END scs8ls_mux2_2

MACRO scs8ls_mux2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.35 0.835 1.78 ;
        RECT 0.665 1.78 0.835 2.05 ;
        RECT 0.665 2.05 1.675 2.155 ;
        RECT 0.665 2.155 3.165 2.22 ;
        RECT 1.505 2.22 3.165 2.325 ;
        RECT 2.995 1.765 3.165 2.155 ;
        RECT 2.995 1.435 3.745 1.765 ;
    END
    ANTENNAGATEAREA 0.738 ;
  END S

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.37 2.755 1.71 ;
        RECT 1.085 1.71 2.77 1.88 ;
        RECT 1.31 0.37 1.64 1.37 ;
        RECT 2.33 0.37 2.755 1.37 ;
        RECT 2.44 1.88 2.77 1.985 ;
    END
    ANTENNADIFFAREA 1.57655 ;
  END X

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.325 1.45 8.175 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.64 1.45 7.075 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A0

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.085 2.495 3.505 2.56 ;
      RECT 1.165 2.56 3.505 2.665 ;
      RECT 3.335 2.105 3.505 2.495 ;
      RECT 3.335 1.935 4.085 2.105 ;
      RECT 3.915 1.765 4.085 1.935 ;
      RECT 3.915 1.435 4.985 1.765 ;
      RECT 0.085 1.15 0.255 1.95 ;
      RECT 0.085 2.56 0.445 2.86 ;
      RECT 0.085 1.95 0.445 2.39 ;
      RECT 0.085 0.47 0.6 1.15 ;
      RECT 0.085 2.39 1.335 2.495 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 1.82 2.835 2.15 3.245 ;
      RECT 3.06 2.835 3.39 3.245 ;
      RECT 4.13 2.775 4.46 3.245 ;
      RECT 5.2 2.775 5.45 3.245 ;
      RECT 0.65 2.73 0.995 3.245 ;
      RECT 8.195 2.2 8.525 2.98 ;
      RECT 6.3 1.95 8.525 2.2 ;
      RECT 8.355 1.03 8.525 1.95 ;
      RECT 8.19 0.425 8.525 1.03 ;
      RECT 5.835 0.255 8.525 0.425 ;
      RECT 7.26 0.425 7.59 0.94 ;
      RECT 6.3 1.78 6.47 1.95 ;
      RECT 5.385 1.45 6.47 1.78 ;
      RECT 5.835 0.425 6.59 0.6 ;
      RECT 7.695 2.54 8.025 2.98 ;
      RECT 5.96 2.37 8.025 2.54 ;
      RECT 5.96 2.265 6.13 2.37 ;
      RECT 4.665 2.095 6.13 2.265 ;
      RECT 4.665 1.935 5.14 2.095 ;
      RECT 5.155 1.265 8.02 1.28 ;
      RECT 3.52 1.11 8.02 1.265 ;
      RECT 3.52 1.095 5.325 1.11 ;
      RECT 7.77 0.595 8.02 1.11 ;
      RECT 3.52 0.575 3.85 1.095 ;
      RECT 0 -0.085 8.64 0.085 ;
      RECT 2.925 0.085 3.255 1.255 ;
      RECT 4.02 0.085 4.49 0.905 ;
      RECT 5.17 0.085 5.575 0.585 ;
      RECT 0.77 0.085 1.1 1.15 ;
      RECT 1.81 0.085 2.14 1.07 ;
      RECT 5.62 2.71 7.115 2.98 ;
      RECT 5.62 2.605 5.79 2.71 ;
      RECT 3.675 2.435 5.79 2.605 ;
      RECT 3.675 2.605 3.925 2.975 ;
      RECT 3.675 2.275 3.925 2.435 ;
      RECT 5.495 0.925 7.09 0.94 ;
      RECT 4.66 0.77 7.09 0.925 ;
      RECT 4.66 0.755 5.665 0.77 ;
      RECT 6.76 0.595 7.09 0.77 ;
      RECT 4.66 0.575 4.99 0.755 ;
    LAYER mcon ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_mux2_4

MACRO scs8ls_mux2i_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.495 0.705 3.225 1.035 ;
        RECT 3.035 1.035 3.225 2.735 ;
    END
    ANTENNADIFFAREA 0.8577 ;
  END Y

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.35 2.865 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395 1.18 3.725 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.55 1.855 ;
    END
    ANTENNAGATEAREA 0.488 ;
  END S

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.08 2.12 1.33 2.98 ;
      RECT 1.08 1.95 2.835 2.12 ;
      RECT 2.505 2.12 2.835 2.735 ;
      RECT 1.08 1.82 1.33 1.95 ;
      RECT 2.06 2.905 3.735 3.075 ;
      RECT 3.405 1.82 3.735 2.905 ;
      RECT 2.06 2.29 2.31 2.905 ;
      RECT 0.555 2.1 0.89 2.98 ;
      RECT 0.72 1.52 0.89 2.1 ;
      RECT 0.72 1.35 2.13 1.52 ;
      RECT 1.8 1.52 2.13 1.68 ;
      RECT 0.72 0.905 0.89 1.35 ;
      RECT 0.545 0.405 0.89 0.905 ;
      RECT 2.105 0.35 3.68 0.52 ;
      RECT 3.395 0.52 3.68 1.01 ;
      RECT 1.105 1.01 2.275 1.18 ;
      RECT 2.105 0.52 2.275 1.01 ;
      RECT 1.105 0.35 1.435 1.01 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 0.115 0.085 0.365 0.905 ;
      RECT 1.605 0.085 1.935 0.84 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 1.53 2.29 1.86 3.245 ;
      RECT 0.105 2.1 0.355 3.245 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_mux2i_1

MACRO scs8ls_mux2i_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535 1.43 3.235 1.775 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.43 4.675 1.84 ;
        RECT 4.35 1.84 5.81 2.01 ;
        RECT 5.48 1.35 5.81 1.84 ;
    END
    ANTENNAGATEAREA 0.804 ;
  END S

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.945 2.845 2.115 ;
        RECT 0.085 2.115 0.445 2.98 ;
        RECT 0.085 1.82 0.445 1.945 ;
        RECT 0.085 1.01 0.255 1.82 ;
        RECT 0.085 0.425 0.45 1.01 ;
        RECT 0.085 0.255 2.91 0.425 ;
        RECT 2.58 0.425 2.91 0.58 ;
    END
    ANTENNADIFFAREA 2.04095 ;
  END Y

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.18 1.315 1.55 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A0

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.685 2.795 2.395 2.955 ;
      RECT 1.685 2.68 3.525 2.795 ;
      RECT 1.685 2.625 5.09 2.68 ;
      RECT 4.76 2.68 5.09 2.98 ;
      RECT 3.355 2.51 5.09 2.625 ;
      RECT 4.76 2.18 5.09 2.51 ;
      RECT 5.795 2.18 6.15 2.86 ;
      RECT 5.98 1.18 6.15 2.18 ;
      RECT 4.91 1.01 6.15 1.18 ;
      RECT 5.795 0.57 6.15 1.01 ;
      RECT 4.91 1.18 5.24 1.67 ;
      RECT 0 3.245 6.24 3.415 ;
      RECT 3.075 2.965 3.47 3.245 ;
      RECT 4.21 2.85 4.555 3.245 ;
      RECT 5.26 2.18 5.59 3.245 ;
      RECT 3.14 0.085 3.47 0.49 ;
      RECT 0 -0.085 6.24 0.085 ;
      RECT 4.21 0.085 4.555 0.49 ;
      RECT 5.285 0.085 5.615 0.84 ;
      RECT 1.74 1.09 4.03 1.26 ;
      RECT 3.65 1 4.03 1.09 ;
      RECT 1.74 0.935 2.07 1.09 ;
      RECT 2.24 0.83 3.25 0.92 ;
      RECT 2.24 0.765 5.115 0.83 ;
      RECT 0.64 0.75 5.115 0.765 ;
      RECT 3.08 0.66 5.115 0.75 ;
      RECT 4.735 0.5 5.115 0.66 ;
      RECT 0.64 0.765 0.97 1.01 ;
      RECT 0.64 0.595 2.41 0.75 ;
      RECT 0.615 2.455 0.945 2.98 ;
      RECT 0.615 2.34 3.185 2.455 ;
      RECT 0.615 2.285 4.005 2.34 ;
      RECT 3.015 2.01 4.005 2.285 ;
    LAYER mcon ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_mux2i_2

MACRO scs8ls_mux2i_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.55 4.245 1.95 ;
        RECT 0.115 1.95 4.245 2.12 ;
        RECT 3.915 1.18 4.085 1.55 ;
        RECT 0.115 2.12 0.365 2.98 ;
        RECT 1.095 2.12 1.265 2.735 ;
        RECT 1.915 2.12 2.245 2.735 ;
        RECT 2.915 2.12 3.245 2.395 ;
        RECT 3.915 2.12 4.245 2.395 ;
        RECT 0.115 1.82 0.365 1.95 ;
        RECT 0.115 1.01 4.085 1.18 ;
        RECT 0.115 1.18 0.365 1.185 ;
        RECT 1.92 0.935 4.085 1.01 ;
        RECT 1.055 0.595 1.225 1.01 ;
        RECT 0.115 0.405 0.365 1.01 ;
        RECT 1.92 0.595 2.25 0.935 ;
    END
    ANTENNADIFFAREA 2.8687 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 1.35 1.885 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.225 1.35 3.235 1.68 ;
        RECT 2.525 1.68 3.235 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A0

  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.08 1.18 9.475 1.54 ;
    END
    ANTENNAGATEAREA 1.479 ;
  END S

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.565 2.905 6.56 3.075 ;
      RECT 5.3 2.73 6.56 2.905 ;
      RECT 0.565 2.29 0.895 2.905 ;
      RECT 1.465 2.29 1.715 2.905 ;
      RECT 4.255 1 6.715 1.17 ;
      RECT 6.385 0.92 6.715 1 ;
      RECT 4.255 0.765 4.425 1 ;
      RECT 2.42 0.595 4.425 0.765 ;
      RECT 7.405 0.84 8.825 1.01 ;
      RECT 7.405 0.75 7.735 0.84 ;
      RECT 8.495 0.39 8.825 0.84 ;
      RECT 4.595 0.66 7.735 0.75 ;
      RECT 4.595 0.75 5.525 0.83 ;
      RECT 5.355 0.58 7.735 0.66 ;
      RECT 4.595 0.425 4.765 0.66 ;
      RECT 7.405 0.39 7.735 0.58 ;
      RECT 0.545 0.255 4.765 0.425 ;
      RECT 0.545 0.425 0.875 0.84 ;
      RECT 1.405 0.425 1.735 0.84 ;
      RECT 2.415 2.565 5.13 2.735 ;
      RECT 4.96 2.56 5.13 2.565 ;
      RECT 4.96 2.39 8.56 2.56 ;
      RECT 7.23 2.56 7.56 2.98 ;
      RECT 8.23 2.56 8.56 2.98 ;
      RECT 2.415 2.29 2.745 2.565 ;
      RECT 3.415 2.29 3.745 2.565 ;
      RECT 9.185 1.88 9.455 2.7 ;
      RECT 6.67 1.71 9.825 1.88 ;
      RECT 9.655 1.01 9.825 1.71 ;
      RECT 9.495 0.39 9.825 1.01 ;
      RECT 6.67 1.67 6.84 1.71 ;
      RECT 5.15 1.34 6.84 1.67 ;
      RECT 0 3.245 10.08 3.415 ;
      RECT 6.73 2.73 7.06 3.245 ;
      RECT 7.73 2.73 8.06 3.245 ;
      RECT 8.76 2.22 9.01 3.245 ;
      RECT 9.635 2.05 9.965 3.245 ;
      RECT 4.475 2.05 9.01 2.22 ;
      RECT 4.475 1.84 6.08 2.05 ;
      RECT 4.935 0.085 5.185 0.49 ;
      RECT 0 -0.085 10.08 0.085 ;
      RECT 5.875 0.085 6.205 0.41 ;
      RECT 6.895 0.085 7.225 0.41 ;
      RECT 7.905 0.085 8.325 0.64 ;
      RECT 8.995 0.085 9.325 1.01 ;
    LAYER mcon ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
  END
END scs8ls_mux2i_4

MACRO scs8ls_mux4_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.08 0.4 9.485 1.18 ;
        RECT 9.245 1.18 9.485 2.56 ;
        RECT 9.22 2.56 9.485 2.89 ;
    END
    ANTENNADIFFAREA 0.5581 ;
  END X

  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.205 1.35 8.535 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END S1

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.99 1.215 1.32 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3 1.215 3.33 2.15 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.5 1.215 3.87 2.15 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.85 1.445 6.18 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A3

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.45 1.215 0.82 1.78 ;
    END
    ANTENNAGATEAREA 0.738 ;
  END S0

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 6.79 2.905 8.52 3.075 ;
      RECT 8.35 2.12 8.52 2.905 ;
      RECT 8.35 1.95 8.915 2.12 ;
      RECT 8.745 1.68 8.915 1.95 ;
      RECT 8.745 1.35 9.075 1.68 ;
      RECT 6.79 1.285 7.12 2.905 ;
      RECT 6.745 1.115 7.12 1.285 ;
      RECT 6.745 0.955 6.925 1.115 ;
      RECT 2.46 0.875 4.75 1.045 ;
      RECT 4.08 1.045 4.41 1.45 ;
      RECT 4.58 1.045 4.75 1.445 ;
      RECT 4.58 1.445 5.34 1.775 ;
      RECT 0.11 0.86 1.7 1.03 ;
      RECT 1.53 1.03 1.7 1.2 ;
      RECT 1.53 0.425 1.7 0.86 ;
      RECT 1.53 1.2 1.86 1.53 ;
      RECT 1.53 0.255 2.63 0.425 ;
      RECT 2.46 0.425 2.63 0.875 ;
      RECT 2.46 1.045 2.79 1.45 ;
      RECT 0.11 1.95 0.555 2.88 ;
      RECT 0.11 1.03 0.28 1.95 ;
      RECT 0.11 0.35 0.445 0.86 ;
      RECT 5.35 2.335 6.62 2.505 ;
      RECT 6.29 2.505 6.62 2.98 ;
      RECT 6.29 1.95 6.62 2.335 ;
      RECT 6.405 0.785 6.575 1.95 ;
      RECT 6.405 0.615 7.355 0.785 ;
      RECT 7.105 0.785 7.355 0.935 ;
      RECT 7.105 0.605 7.355 0.615 ;
      RECT 3.795 2.905 5.55 3.075 ;
      RECT 3.795 2.505 4.02 2.905 ;
      RECT 5.35 2.505 5.55 2.905 ;
      RECT 2.03 2.335 4.02 2.505 ;
      RECT 2.03 2.505 2.55 2.725 ;
      RECT 2.03 1.685 2.55 2.335 ;
      RECT 2.03 1.03 2.2 1.685 ;
      RECT 1.875 0.595 2.2 1.03 ;
      RECT 4.92 1.105 6.235 1.275 ;
      RECT 5.985 0.445 6.235 1.105 ;
      RECT 5.985 0.435 6.485 0.445 ;
      RECT 5.985 0.265 7.695 0.435 ;
      RECT 7.525 0.435 7.695 1.105 ;
      RECT 7.29 1.105 7.695 1.275 ;
      RECT 7.29 1.275 7.46 1.945 ;
      RECT 7.29 1.945 7.62 2.735 ;
      RECT 4.305 2.165 5.165 2.735 ;
      RECT 4.305 1.995 5.68 2.165 ;
      RECT 5.51 1.275 5.68 1.995 ;
      RECT 4.92 0.705 5.09 1.105 ;
      RECT 4.21 0.375 5.09 0.705 ;
      RECT 7.865 0.5 8.41 1.18 ;
      RECT 7.85 1.95 8.18 2.735 ;
      RECT 7.85 1.775 8.035 1.95 ;
      RECT 7.63 1.445 8.035 1.775 ;
      RECT 7.865 1.18 8.035 1.445 ;
      RECT 0 -0.085 9.6 0.085 ;
      RECT 0.7 0.085 1.09 0.68 ;
      RECT 3.125 0.085 3.715 0.68 ;
      RECT 5.26 0.085 5.59 0.935 ;
      RECT 8.58 0.085 8.91 1.18 ;
      RECT 0 3.245 9.6 3.415 ;
      RECT 3.265 2.675 3.595 3.245 ;
      RECT 5.73 2.675 6.06 3.245 ;
      RECT 8.69 2.29 9.02 3.245 ;
      RECT 0.725 1.95 1.055 3.245 ;
    LAYER mcon ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
  END
END scs8ls_mux4_1

MACRO scs8ls_dlxtn_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805 1.15 8.035 1.82 ;
        RECT 6.315 1.82 8.035 1.99 ;
        RECT 6.265 0.98 8.035 1.15 ;
        RECT 7.315 1.99 8.035 2.15 ;
        RECT 6.315 1.99 6.645 2.98 ;
        RECT 6.265 0.35 6.615 0.98 ;
        RECT 7.295 0.35 7.545 0.98 ;
        RECT 7.315 2.15 7.545 2.98 ;
    END
    ANTENNADIFFAREA 1.2703 ;
  END Q

  PIN GATEN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.985 1.5 1.315 1.83 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END GATEN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.3 0.455 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.36 2.06 3.88 2.735 ;
      RECT 3.71 1.055 3.88 2.06 ;
      RECT 3.655 0.725 4.72 1.055 ;
      RECT 4.55 1.055 4.72 1.32 ;
      RECT 4.55 1.32 5.49 1.65 ;
      RECT 1.825 1.94 2.225 2.22 ;
      RECT 2.055 1.89 2.225 1.94 ;
      RECT 2.055 1.72 3.54 1.89 ;
      RECT 3.21 1.47 3.54 1.72 ;
      RECT 2.055 0.595 2.305 1.72 ;
      RECT 3.315 0.505 3.485 1.47 ;
      RECT 3.315 0.255 4.445 0.505 ;
      RECT 5.66 1.32 7.49 1.65 ;
      RECT 5.315 2.305 5.645 2.98 ;
      RECT 4.39 1.99 5.645 2.305 ;
      RECT 4.39 1.975 5.83 1.99 ;
      RECT 5.315 1.82 5.83 1.975 ;
      RECT 5.66 1.65 5.83 1.82 ;
      RECT 5.66 1.15 5.83 1.32 ;
      RECT 5.32 0.98 5.83 1.15 ;
      RECT 5.32 0.375 5.57 0.98 ;
      RECT 1.135 2.56 1.655 2.98 ;
      RECT 1.135 2.39 3.16 2.56 ;
      RECT 2.99 2.56 3.16 2.905 ;
      RECT 1.135 2.1 1.655 2.39 ;
      RECT 2.99 2.905 4.22 3.075 ;
      RECT 1.485 1.77 1.655 2.1 ;
      RECT 4.05 1.735 4.22 2.905 ;
      RECT 1.485 1.33 1.885 1.77 ;
      RECT 4.05 1.405 4.38 1.735 ;
      RECT 1.135 1 1.885 1.33 ;
      RECT 1.485 0.76 1.885 1 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 7.715 0.085 8.045 0.81 ;
      RECT 0.625 0.085 0.955 0.49 ;
      RECT 2.815 0.085 3.145 1.05 ;
      RECT 4.89 0.085 5.14 1.055 ;
      RECT 5.75 0.085 6.08 0.81 ;
      RECT 6.785 0.085 7.115 0.81 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 7.715 2.32 8.045 3.245 ;
      RECT 2.36 2.73 2.82 3.245 ;
      RECT 4.39 2.59 5.145 3.245 ;
      RECT 0.635 2.29 0.965 3.245 ;
      RECT 5.815 2.16 6.145 3.245 ;
      RECT 6.815 2.16 7.145 3.245 ;
      RECT 0.115 0.66 1.315 0.83 ;
      RECT 1.145 0.425 1.315 0.66 ;
      RECT 1.145 0.255 2.645 0.425 ;
      RECT 2.475 0.425 2.645 1.22 ;
      RECT 2.475 1.22 3 1.55 ;
      RECT 0.135 2.12 0.465 2.98 ;
      RECT 0.135 1.95 0.795 2.12 ;
      RECT 0.625 1.13 0.795 1.95 ;
      RECT 0.115 0.83 0.795 1.13 ;
      RECT 0.115 0.555 0.445 0.66 ;
    LAYER mcon ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_dlxtn_4

MACRO scs8ls_dlxtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.35 6.715 1.78 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END GATE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.23 1.82 7.595 2.98 ;
        RECT 7.425 1.15 7.595 1.82 ;
        RECT 7.235 0.39 7.595 1.15 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.595 1.85 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.125 2.785 1.455 2.98 ;
      RECT 1.125 2.735 2.97 2.785 ;
      RECT 2.165 2.785 2.97 2.985 ;
      RECT 1.125 2.615 2.335 2.735 ;
      RECT 1.125 1.94 1.455 2.615 ;
      RECT 1.335 1.355 2.345 1.525 ;
      RECT 1.335 0.93 1.505 1.355 ;
      RECT 2.175 0.925 2.345 1.355 ;
      RECT 1.175 0.405 1.505 0.93 ;
      RECT 2.175 0.765 2.845 0.925 ;
      RECT 2.175 0.755 3.895 0.765 ;
      RECT 2.675 0.595 3.895 0.755 ;
      RECT 3.14 2.845 4.04 3.015 ;
      RECT 3.14 2.565 3.31 2.845 ;
      RECT 2.505 2.445 3.31 2.565 ;
      RECT 2.08 2.395 3.31 2.445 ;
      RECT 2.08 2.275 2.675 2.395 ;
      RECT 2.08 1.94 2.33 2.275 ;
      RECT 6.895 1.32 7.255 1.65 ;
      RECT 4.565 0.58 7.065 0.75 ;
      RECT 6.895 0.75 7.065 1.32 ;
      RECT 4.27 1.665 4.815 1.995 ;
      RECT 4.565 0.75 4.815 1.665 ;
      RECT 4.565 0.425 4.815 0.58 ;
      RECT 2.175 0.255 4.815 0.425 ;
      RECT 2.175 0.425 2.505 0.585 ;
      RECT 0.645 2.1 0.945 2.98 ;
      RECT 0.775 1.77 0.945 2.1 ;
      RECT 0.775 1.1 1.165 1.77 ;
      RECT 0.775 1.01 0.945 1.1 ;
      RECT 0.615 0.42 0.945 1.01 ;
      RECT 3.93 2.165 5.625 2.335 ;
      RECT 3.93 1.545 4.1 2.165 ;
      RECT 5.375 1.17 5.625 2.165 ;
      RECT 3.525 1.275 4.1 1.545 ;
      RECT 5.375 0.92 5.835 1.17 ;
      RECT 2.845 2.105 3.42 2.225 ;
      RECT 2.515 2.055 3.42 2.105 ;
      RECT 2.515 1.935 3.015 2.055 ;
      RECT 2.515 1.265 2.685 1.935 ;
      RECT 2.515 1.105 3.355 1.265 ;
      RECT 2.515 1.095 4.395 1.105 ;
      RECT 3.015 0.935 4.395 1.095 ;
      RECT 4.065 0.775 4.395 0.935 ;
      RECT 5.34 2.675 6.525 2.7 ;
      RECT 3.59 2.505 6.525 2.675 ;
      RECT 5.845 1.95 6.525 2.505 ;
      RECT 6.005 0.92 6.41 1.17 ;
      RECT 3.59 1.885 3.76 2.505 ;
      RECT 5.845 1.35 6.175 1.95 ;
      RECT 3.185 1.765 3.76 1.885 ;
      RECT 6.005 1.17 6.175 1.35 ;
      RECT 2.855 1.715 3.76 1.765 ;
      RECT 2.855 1.435 3.355 1.715 ;
      RECT 0 -0.085 7.68 0.085 ;
      RECT 0.115 0.085 0.445 1.01 ;
      RECT 1.675 0.085 2.005 1.185 ;
      RECT 4.995 0.085 5.325 0.41 ;
      RECT 6.59 0.085 7.055 0.41 ;
      RECT 0 3.245 7.68 3.415 ;
      RECT 1.66 2.955 1.995 3.245 ;
      RECT 4.84 2.845 5.17 3.245 ;
      RECT 0.115 2.1 0.445 3.245 ;
      RECT 6.73 1.95 7.06 3.245 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
  END
END scs8ls_dlxtp_1

MACRO scs8ls_dlygate4sd1_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.45 1.12 3.74 1.815 ;
        RECT 3.325 1.815 3.74 3.06 ;
        RECT 3.325 0.355 3.74 1.12 ;
    END
    ANTENNADIFFAREA 0.5097 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.19 0.73 1.86 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END A

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 0.585 0.085 0.915 0.65 ;
      RECT 2.825 0.085 3.155 0.87 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 0.575 2.38 0.905 3.245 ;
      RECT 2.825 2.165 3.155 3.245 ;
      RECT 1.985 1.995 2.345 2.19 ;
      RECT 1.985 1.825 3.155 1.995 ;
      RECT 2.91 1.625 3.155 1.825 ;
      RECT 2.91 1.295 3.28 1.625 ;
      RECT 2.91 1.21 3.155 1.295 ;
      RECT 1.985 1.04 3.155 1.21 ;
      RECT 1.985 0.71 2.345 1.04 ;
      RECT 1.415 2.395 1.72 2.725 ;
      RECT 1.475 1.61 1.72 2.395 ;
      RECT 1.475 1.38 2.74 1.61 ;
      RECT 1.475 0.635 1.72 1.38 ;
      RECT 1.415 0.305 1.72 0.635 ;
      RECT 0.095 2.205 0.4 2.725 ;
      RECT 0.095 2.03 1.305 2.205 ;
      RECT 0.975 1.02 1.305 2.03 ;
      RECT 0.095 0.82 1.305 1.02 ;
      RECT 0.095 0.305 0.41 0.82 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_dlygate4sd1_1

MACRO scs8ls_dlygate4sd2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.45 1.12 3.74 1.815 ;
        RECT 3.325 1.815 3.74 3.06 ;
        RECT 3.325 0.355 3.74 1.12 ;
    END
    ANTENNADIFFAREA 0.5097 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.19 0.73 1.86 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END A

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 0.585 0.085 0.915 0.65 ;
      RECT 2.825 0.085 3.155 0.87 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 0.575 2.38 0.905 3.245 ;
      RECT 2.825 2.165 3.155 3.245 ;
      RECT 1.985 1.995 2.345 2.19 ;
      RECT 1.985 1.825 3.155 1.995 ;
      RECT 2.91 1.625 3.155 1.825 ;
      RECT 2.91 1.295 3.28 1.625 ;
      RECT 2.91 1.21 3.155 1.295 ;
      RECT 1.985 1.04 3.155 1.21 ;
      RECT 1.985 0.71 2.345 1.04 ;
      RECT 1.415 2.395 1.72 2.725 ;
      RECT 1.475 1.61 1.72 2.395 ;
      RECT 1.475 1.38 2.74 1.61 ;
      RECT 1.475 0.635 1.72 1.38 ;
      RECT 1.415 0.305 1.72 0.635 ;
      RECT 0.095 2.205 0.4 2.725 ;
      RECT 0.095 2.03 1.305 2.205 ;
      RECT 0.975 1.02 1.305 2.03 ;
      RECT 0.095 0.82 1.305 1.02 ;
      RECT 0.095 0.305 0.41 0.82 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_dlygate4sd2_1

MACRO scs8ls_dlygate4sd3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.45 1.12 3.74 1.815 ;
        RECT 3.325 1.815 3.74 3.06 ;
        RECT 3.325 0.355 3.74 1.12 ;
    END
    ANTENNADIFFAREA 0.5097 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.19 0.73 1.86 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END A

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 0.585 0.085 0.915 0.65 ;
      RECT 2.825 0.085 3.155 0.87 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 0.575 2.38 0.905 3.245 ;
      RECT 2.825 2.165 3.155 3.245 ;
      RECT 1.985 1.995 2.345 2.19 ;
      RECT 1.985 1.825 3.155 1.995 ;
      RECT 2.91 1.625 3.155 1.825 ;
      RECT 2.91 1.295 3.28 1.625 ;
      RECT 2.91 1.21 3.155 1.295 ;
      RECT 1.985 1.04 3.155 1.21 ;
      RECT 1.985 0.71 2.345 1.04 ;
      RECT 1.415 2.395 1.72 2.725 ;
      RECT 1.475 1.61 1.72 2.395 ;
      RECT 1.475 1.38 2.74 1.61 ;
      RECT 1.475 0.635 1.72 1.38 ;
      RECT 1.415 0.305 1.72 0.635 ;
      RECT 0.095 2.205 0.4 2.725 ;
      RECT 0.095 2.03 1.305 2.205 ;
      RECT 0.975 1.02 1.305 2.03 ;
      RECT 0.095 0.82 1.305 1.02 ;
      RECT 0.095 0.305 0.41 0.82 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_dlygate4sd3_1

MACRO scs8ls_dlymetal6s2s_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.355 0.555 1.765 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.965 2.32 4.21 2.49 ;
        RECT 0.965 1.92 1.345 2.32 ;
    END
    ANTENNADIFFAREA 0.5041 ;
    ANTENNAGATEAREA 0.126 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.28 LAYER met1 ;
  END X

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 3.845 1.92 4.225 2.15 ;
      RECT 2.405 1.92 2.785 2.15 ;
    LAYER li1 ;
      RECT 0.1 2.14 0.43 2.225 ;
      RECT 0.1 1.935 0.895 2.14 ;
      RECT 0.725 1.605 0.895 1.935 ;
      RECT 0.725 1.275 1.04 1.605 ;
      RECT 0.725 1.145 0.895 1.275 ;
      RECT 0.1 0.975 0.895 1.145 ;
      RECT 0.1 0.7 0.395 0.975 ;
      RECT 1.065 1.835 1.38 3.075 ;
      RECT 1.21 1.605 1.38 1.835 ;
      RECT 1.21 1.315 1.995 1.605 ;
      RECT 1.21 1.075 1.38 1.315 ;
      RECT 1.09 0.255 1.38 1.075 ;
      RECT 1.55 2.14 1.87 2.225 ;
      RECT 1.55 1.895 2.335 2.14 ;
      RECT 2.165 1.605 2.335 1.895 ;
      RECT 2.165 1.275 2.525 1.605 ;
      RECT 2.165 1.145 2.335 1.275 ;
      RECT 1.55 0.975 2.335 1.145 ;
      RECT 1.55 0.7 1.835 0.975 ;
      RECT 2.565 2.16 2.865 3.075 ;
      RECT 2.505 1.835 2.865 2.16 ;
      RECT 2.695 1.605 2.865 1.835 ;
      RECT 2.695 1.315 3.435 1.605 ;
      RECT 2.695 1.075 2.865 1.315 ;
      RECT 2.53 0.255 2.865 1.075 ;
      RECT 3.07 2.14 3.4 2.225 ;
      RECT 3.07 1.895 3.805 2.14 ;
      RECT 3.605 1.605 3.805 1.895 ;
      RECT 3.605 1.275 4.01 1.605 ;
      RECT 3.605 1.145 3.775 1.275 ;
      RECT 3.06 0.975 3.775 1.145 ;
      RECT 3.06 0.7 3.275 0.975 ;
      RECT 4.05 2.16 4.35 3.075 ;
      RECT 3.975 1.835 4.35 2.16 ;
      RECT 4.18 1.075 4.35 1.835 ;
      RECT 3.97 0.255 4.35 1.075 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 0.59 2.31 0.885 3.245 ;
      RECT 2.1 2.31 2.395 3.245 ;
      RECT 3.585 2.31 3.88 3.245 ;
      RECT 0.59 0.085 0.92 0.805 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 2.03 0.085 2.36 0.805 ;
      RECT 3.47 0.085 3.8 0.805 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 1.115 1.95 1.285 2.12 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 2.555 1.95 2.725 2.12 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.995 1.95 4.165 2.12 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
  END
END scs8ls_dlymetal6s2s_1

MACRO scs8ls_dlymetal6s4s_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.355 0.555 1.765 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.965 2.32 4.21 2.49 ;
        RECT 2.405 1.92 2.785 2.32 ;
    END
    ANTENNADIFFAREA 0.5041 ;
    ANTENNAGATEAREA 0.126 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.28 LAYER met1 ;
  END X

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 3.845 1.92 4.225 2.15 ;
      RECT 0.965 1.92 1.345 2.15 ;
    LAYER li1 ;
      RECT 0.1 2.14 0.43 2.225 ;
      RECT 0.1 1.935 0.895 2.14 ;
      RECT 0.725 1.605 0.895 1.935 ;
      RECT 0.725 1.275 1.04 1.605 ;
      RECT 0.725 1.145 0.895 1.275 ;
      RECT 0.1 0.975 0.895 1.145 ;
      RECT 0.1 0.7 0.395 0.975 ;
      RECT 1.065 1.835 1.38 3.075 ;
      RECT 1.21 1.605 1.38 1.835 ;
      RECT 1.21 1.315 1.995 1.605 ;
      RECT 1.21 1.075 1.38 1.315 ;
      RECT 1.09 0.255 1.38 1.075 ;
      RECT 1.55 2.14 1.87 2.225 ;
      RECT 1.55 1.895 2.335 2.14 ;
      RECT 2.165 1.605 2.335 1.895 ;
      RECT 2.165 1.275 2.525 1.605 ;
      RECT 2.165 1.145 2.335 1.275 ;
      RECT 1.55 0.975 2.335 1.145 ;
      RECT 1.55 0.7 1.835 0.975 ;
      RECT 2.565 2.16 2.865 3.075 ;
      RECT 2.505 1.835 2.865 2.16 ;
      RECT 2.695 1.605 2.865 1.835 ;
      RECT 2.695 1.315 3.435 1.605 ;
      RECT 2.695 1.075 2.865 1.315 ;
      RECT 2.53 0.255 2.865 1.075 ;
      RECT 3.07 2.14 3.4 2.225 ;
      RECT 3.07 1.895 3.805 2.14 ;
      RECT 3.605 1.605 3.805 1.895 ;
      RECT 3.605 1.275 4.01 1.605 ;
      RECT 3.605 1.145 3.775 1.275 ;
      RECT 3.06 0.975 3.775 1.145 ;
      RECT 3.06 0.7 3.275 0.975 ;
      RECT 4.05 2.16 4.35 3.075 ;
      RECT 3.975 1.835 4.35 2.16 ;
      RECT 4.18 1.075 4.35 1.835 ;
      RECT 3.97 0.255 4.35 1.075 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 0.59 2.31 0.885 3.245 ;
      RECT 2.1 2.31 2.395 3.245 ;
      RECT 3.585 2.31 3.88 3.245 ;
      RECT 0.59 0.085 0.92 0.805 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 2.03 0.085 2.36 0.805 ;
      RECT 3.47 0.085 3.8 0.805 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 1.115 1.95 1.285 2.12 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 2.555 1.95 2.725 2.12 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.995 1.95 4.165 2.12 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
  END
END scs8ls_dlymetal6s4s_1

MACRO scs8ls_dlymetal6s6s_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.355 0.555 1.765 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3.845 1.92 4.225 2.32 ;
        RECT 0.965 2.32 4.225 2.49 ;
    END
    ANTENNADIFFAREA 0.5041 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2905 LAYER met1 ;
  END X

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 0.965 1.92 1.345 2.15 ;
      RECT 2.405 1.92 2.785 2.15 ;
    LAYER li1 ;
      RECT 0.1 2.14 0.43 2.225 ;
      RECT 0.1 1.935 0.895 2.14 ;
      RECT 0.725 1.605 0.895 1.935 ;
      RECT 0.725 1.275 1.04 1.605 ;
      RECT 0.725 1.145 0.895 1.275 ;
      RECT 0.1 0.975 0.895 1.145 ;
      RECT 0.1 0.7 0.395 0.975 ;
      RECT 1.065 1.835 1.38 3.075 ;
      RECT 1.21 1.605 1.38 1.835 ;
      RECT 1.21 1.315 1.995 1.605 ;
      RECT 1.21 1.075 1.38 1.315 ;
      RECT 1.09 0.255 1.38 1.075 ;
      RECT 1.55 2.14 1.87 2.225 ;
      RECT 1.55 1.895 2.335 2.14 ;
      RECT 2.165 1.605 2.335 1.895 ;
      RECT 2.165 1.275 2.525 1.605 ;
      RECT 2.165 1.145 2.335 1.275 ;
      RECT 1.55 0.975 2.335 1.145 ;
      RECT 1.55 0.7 1.835 0.975 ;
      RECT 2.565 2.16 2.865 3.075 ;
      RECT 2.505 1.835 2.865 2.16 ;
      RECT 2.695 1.605 2.865 1.835 ;
      RECT 2.695 1.315 3.435 1.605 ;
      RECT 2.695 1.075 2.865 1.315 ;
      RECT 2.53 0.255 2.865 1.075 ;
      RECT 3.07 2.14 3.4 2.225 ;
      RECT 3.07 1.895 3.805 2.14 ;
      RECT 3.605 1.605 3.805 1.895 ;
      RECT 3.605 1.275 4.01 1.605 ;
      RECT 3.605 1.145 3.775 1.275 ;
      RECT 3.06 0.975 3.775 1.145 ;
      RECT 3.06 0.7 3.275 0.975 ;
      RECT 4.05 2.16 4.35 3.075 ;
      RECT 3.975 1.835 4.35 2.16 ;
      RECT 4.18 1.075 4.35 1.835 ;
      RECT 3.97 0.255 4.35 1.075 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 0.59 2.31 0.885 3.245 ;
      RECT 2.1 2.31 2.395 3.245 ;
      RECT 3.585 2.31 3.88 3.245 ;
      RECT 0.59 0.085 0.92 0.805 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 2.03 0.085 2.36 0.805 ;
      RECT 3.47 0.085 3.8 0.805 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 1.115 1.95 1.285 2.12 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 2.555 1.95 2.725 2.12 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.995 1.95 4.165 2.12 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
  END
END scs8ls_dlymetal6s6s_1

MACRO scs8ls_ebufn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.5 0.835 1.83 ;
        RECT 0.665 1.83 0.835 2.42 ;
        RECT 0.665 2.42 2.195 2.59 ;
        RECT 1.865 2.59 2.195 3.01 ;
        RECT 1.865 2.34 2.195 2.42 ;
    END
    ANTENNAGATEAREA 0.377 ;
  END TEB

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.21 0.35 3.755 1.13 ;
        RECT 3.585 1.13 3.755 1.82 ;
        RECT 3.235 1.82 3.755 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END Z

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.5 1.795 1.83 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.46 1.32 3.415 1.65 ;
      RECT 1.185 2.17 1.695 2.25 ;
      RECT 1.185 2 2.135 2.17 ;
      RECT 1.965 1.88 2.135 2 ;
      RECT 1.965 1.71 3.065 1.88 ;
      RECT 2.46 1.65 3.065 1.71 ;
      RECT 2.46 0.98 2.66 1.32 ;
      RECT 1.155 0.81 2.66 0.98 ;
      RECT 1.155 0.455 1.45 0.81 ;
      RECT 0.085 1.15 2.2 1.32 ;
      RECT 1.87 1.32 2.2 1.34 ;
      RECT 0.085 1.32 0.255 2 ;
      RECT 0.085 2 0.445 2.88 ;
      RECT 0.085 0.455 0.53 1.15 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 2.365 2.05 2.695 3.245 ;
      RECT 0.65 2.76 0.98 3.245 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 0.7 0.085 0.985 0.85 ;
      RECT 2.39 0.085 2.72 0.64 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_ebufn_1

MACRO scs8ls_ebufn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.35 3.865 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A

  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.965 1.18 3.295 1.65 ;
    END
    ANTENNAGATEAREA 0.582 ;
  END TEB

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.645 1.97 1.795 2.15 ;
        RECT 0.535 1.8 1.795 1.97 ;
        RECT 0.645 2.15 0.975 2.735 ;
        RECT 0.535 1.13 0.705 1.8 ;
        RECT 0.535 0.615 0.875 1.13 ;
    END
    ANTENNADIFFAREA 0.5992 ;
  END Z

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.115 0.255 1.375 0.425 ;
      RECT 1.045 0.425 1.375 0.96 ;
      RECT 1.045 0.96 2.225 1.13 ;
      RECT 1.975 0.35 2.225 0.96 ;
      RECT 0.115 0.425 0.365 1.13 ;
      RECT 0.145 2.905 1.475 3.075 ;
      RECT 1.145 2.75 1.475 2.905 ;
      RECT 1.145 2.58 2.545 2.75 ;
      RECT 2.215 2.75 2.545 2.98 ;
      RECT 1.145 2.32 1.475 2.58 ;
      RECT 0.145 2.14 0.475 2.905 ;
      RECT 2.395 1.82 3.105 2.07 ;
      RECT 2.395 0.325 3.17 1.01 ;
      RECT 2.395 1.01 2.725 1.82 ;
      RECT 3.875 2.41 4.205 2.86 ;
      RECT 1.965 2.24 4.205 2.41 ;
      RECT 3.875 1.95 4.205 2.24 ;
      RECT 4.035 1.03 4.205 1.95 ;
      RECT 3.84 0.35 4.205 1.03 ;
      RECT 1.965 1.63 2.135 2.24 ;
      RECT 0.875 1.3 2.135 1.63 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 1.68 2.92 2.01 3.245 ;
      RECT 3.225 2.61 3.705 3.245 ;
      RECT 1.545 0.085 1.795 0.79 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 3.34 0.085 3.67 1.01 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_ebufn_2

MACRO scs8ls_ebufn_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.3 0.805 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.975 1.18 1.285 1.55 ;
    END
    ANTENNAGATEAREA 0.951 ;
  END TEB

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.87 1.99 5.205 2.735 ;
        RECT 3.97 1.82 5.205 1.99 ;
        RECT 3.97 1.99 4.3 2.735 ;
        RECT 5.035 1.15 5.205 1.82 ;
        RECT 4.015 0.98 5.205 1.15 ;
        RECT 4.015 0.595 4.345 0.98 ;
        RECT 4.875 0.595 5.205 0.98 ;
    END
    ANTENNADIFFAREA 1.1012 ;
  END Z

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.585 0.255 5.655 0.425 ;
      RECT 5.405 0.425 5.655 1.13 ;
      RECT 1.945 1.15 2.975 1.31 ;
      RECT 1.945 1.14 3.835 1.15 ;
      RECT 2.805 0.98 3.835 1.14 ;
      RECT 1.945 0.35 2.115 1.14 ;
      RECT 3.585 0.425 3.835 0.98 ;
      RECT 2.805 0.35 2.975 0.98 ;
      RECT 4.525 0.425 4.695 0.81 ;
      RECT 3.52 2.905 5.65 3.075 ;
      RECT 5.4 1.82 5.65 2.905 ;
      RECT 3.52 1.99 3.77 2.905 ;
      RECT 2.7 1.82 3.77 1.99 ;
      RECT 2.7 1.99 2.87 2.4 ;
      RECT 1.8 2.4 2.87 2.57 ;
      RECT 1.8 2.57 1.97 2.82 ;
      RECT 2.7 2.57 2.87 2.98 ;
      RECT 4.47 2.16 4.7 2.905 ;
      RECT 2.36 1.48 4.83 1.65 ;
      RECT 3.82 1.32 4.83 1.48 ;
      RECT 0.085 2.39 1.63 2.56 ;
      RECT 1.46 2.23 1.63 2.39 ;
      RECT 1.46 2.06 2.53 2.23 ;
      RECT 2.36 1.65 2.53 2.06 ;
      RECT 0.085 2.56 0.365 2.98 ;
      RECT 0.085 1.95 0.365 2.39 ;
      RECT 0.085 1.13 0.255 1.95 ;
      RECT 0.085 0.35 0.405 1.13 ;
      RECT 1.04 1.89 1.29 2.22 ;
      RECT 1.04 1.72 1.775 1.89 ;
      RECT 1.455 1.01 1.775 1.72 ;
      RECT 1.095 0.3 1.775 1.01 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 2.17 2.74 2.5 3.245 ;
      RECT 0.565 2.73 0.92 3.245 ;
      RECT 3.07 2.16 3.32 3.245 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 0.585 0.085 0.915 1.01 ;
      RECT 2.295 0.085 2.625 0.97 ;
      RECT 3.155 0.085 3.405 0.81 ;
    LAYER mcon ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_ebufn_4

MACRO scs8ls_ebufn_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 0.595 0.875 0.98 ;
        RECT 0.545 0.98 3.76 1.15 ;
        RECT 0.545 1.15 0.835 1.82 ;
        RECT 1.43 0.595 1.76 0.98 ;
        RECT 2.43 0.595 2.76 0.98 ;
        RECT 3.43 0.595 3.76 0.98 ;
        RECT 0.545 1.82 3.7 1.99 ;
        RECT 0.545 1.99 0.9 2.735 ;
        RECT 1.52 1.99 1.85 2.735 ;
        RECT 2.42 1.99 2.75 2.735 ;
        RECT 3.37 1.99 3.7 2.735 ;
    END
    ANTENNADIFFAREA 2.3605 ;
  END Z

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.645 1.18 9.975 1.55 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A

  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.265 1.18 9.475 1.55 ;
    END
    ANTENNAGATEAREA 1.623 ;
  END TEB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 4.72 1.31 7.55 1.47 ;
      RECT 3.94 1.3 7.55 1.31 ;
      RECT 3.94 1.14 5.05 1.3 ;
      RECT 5.58 0.35 5.83 1.3 ;
      RECT 6.44 0.35 6.69 1.3 ;
      RECT 7.3 0.35 7.55 1.3 ;
      RECT 3.94 0.425 4.11 1.14 ;
      RECT 4.8 0.35 5.05 1.14 ;
      RECT 0.115 0.255 4.11 0.425 ;
      RECT 0.115 0.425 0.365 1.13 ;
      RECT 1.055 0.425 1.225 0.81 ;
      RECT 1.93 0.425 2.26 0.81 ;
      RECT 2.93 0.425 3.26 0.81 ;
      RECT 0.12 2.905 4.2 3.075 ;
      RECT 3.87 2.56 4.2 2.905 ;
      RECT 3.87 2.39 7.2 2.56 ;
      RECT 4.87 2.56 5.2 2.98 ;
      RECT 5.87 2.56 6.2 2.98 ;
      RECT 6.87 2.56 8.27 2.73 ;
      RECT 6.87 2.73 7.2 2.98 ;
      RECT 7.94 2.73 8.27 2.98 ;
      RECT 0.12 1.82 0.37 2.905 ;
      RECT 1.085 2.16 1.35 2.905 ;
      RECT 2.05 2.16 2.22 2.905 ;
      RECT 2.92 2.16 3.19 2.905 ;
      RECT 9.665 2.39 9.945 2.98 ;
      RECT 7.585 2.22 9.945 2.39 ;
      RECT 9.665 1.89 9.945 2.22 ;
      RECT 9.665 1.72 10.315 1.89 ;
      RECT 10.145 1.01 10.315 1.72 ;
      RECT 9.68 0.84 10.315 1.01 ;
      RECT 9.68 0.34 9.93 0.84 ;
      RECT 3.87 2.05 7.755 2.22 ;
      RECT 3.87 1.65 4.04 2.05 ;
      RECT 1.035 1.48 4.04 1.65 ;
      RECT 1.035 1.32 3.655 1.48 ;
      RECT 7.925 1.8 9.045 2.05 ;
      RECT 7.925 0.67 9.15 1.01 ;
      RECT 7.72 0.34 9.15 0.67 ;
      RECT 7.925 1.01 8.095 1.8 ;
      RECT 0 3.245 10.56 3.415 ;
      RECT 7.405 2.9 7.735 3.245 ;
      RECT 4.37 2.73 4.7 3.245 ;
      RECT 5.37 2.73 5.7 3.245 ;
      RECT 6.37 2.73 6.7 3.245 ;
      RECT 9.165 2.56 9.495 3.245 ;
      RECT 10.115 2.06 10.445 3.245 ;
      RECT 4.29 0.085 4.62 0.97 ;
      RECT 0 -0.085 10.56 0.085 ;
      RECT 5.23 0.085 5.4 1.13 ;
      RECT 6.01 0.085 6.26 1.13 ;
      RECT 6.87 0.085 7.12 1.13 ;
      RECT 9.33 0.085 9.5 1.01 ;
      RECT 10.11 0.085 10.445 0.6 ;
    LAYER mcon ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
  END
END scs8ls_ebufn_8

MACRO scs8ls_edfxbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 14.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.955 0.37 14.315 1.15 ;
        RECT 14.145 1.15 14.315 1.82 ;
        RECT 13.99 1.82 14.315 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END QN

  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.45 1.905 1.78 ;
    END
    ANTENNAGATEAREA 0.285 ;
  END DE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.98 0.835 1.99 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.925 1.82 13.34 2.98 ;
        RECT 12.925 1 13.095 1.82 ;
        RECT 12.765 0.62 13.095 1 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.715 1.18 4.385 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 12.155 1.58 12.325 1.75 ;
      RECT 3.035 1.58 3.205 1.75 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
    LAYER met1 ;
      RECT 2.975 1.735 3.265 1.78 ;
      RECT 2.975 1.595 12.385 1.735 ;
      RECT 12.095 1.735 12.385 1.78 ;
      RECT 2.975 1.55 3.265 1.595 ;
      RECT 12.095 1.55 12.385 1.595 ;
    LAYER li1 ;
      RECT 8.195 2.755 9.405 2.925 ;
      RECT 8.195 2.715 8.365 2.755 ;
      RECT 9.235 1.79 9.405 2.755 ;
      RECT 7.15 2.545 8.365 2.715 ;
      RECT 9.235 1.62 10.625 1.79 ;
      RECT 7.15 2.38 7.32 2.545 ;
      RECT 10.295 1.46 10.625 1.62 ;
      RECT 6.89 2.08 7.32 2.38 ;
      RECT 1.715 2.12 1.885 2.735 ;
      RECT 1.005 1.95 2.665 2.12 ;
      RECT 2.335 0.98 2.665 1.95 ;
      RECT 1.005 1.11 2 1.28 ;
      RECT 1.65 0.48 2 1.11 ;
      RECT 1.005 1.28 1.335 1.95 ;
      RECT 10.445 2.155 10.775 2.98 ;
      RECT 10.445 1.985 11.445 2.155 ;
      RECT 11.275 1.485 11.445 1.985 ;
      RECT 11.275 1.155 11.985 1.485 ;
      RECT 11.275 0.95 11.445 1.155 ;
      RECT 9.54 0.62 11.445 0.95 ;
      RECT 8.7 2.375 9.03 2.585 ;
      RECT 8.23 2.125 9.03 2.375 ;
      RECT 8.7 1.475 9.03 2.125 ;
      RECT 7.205 1.305 9.03 1.475 ;
      RECT 7.205 1.475 7.535 1.57 ;
      RECT 7.98 0.595 8.15 1.305 ;
      RECT 5.955 2.14 6.355 2.38 ;
      RECT 5.555 1.97 6.355 2.14 ;
      RECT 5.555 1.81 6.125 1.97 ;
      RECT 5.955 0.425 6.125 1.81 ;
      RECT 5.095 0.255 6.885 0.425 ;
      RECT 5.095 0.425 5.345 1.13 ;
      RECT 6.635 0.425 6.885 0.965 ;
      RECT 6.635 0.965 7.81 1.135 ;
      RECT 6.635 1.135 6.885 1.345 ;
      RECT 7.64 0.425 7.81 0.965 ;
      RECT 7.64 0.255 8.49 0.425 ;
      RECT 8.32 0.425 8.49 0.965 ;
      RECT 8.32 0.965 9.37 1.12 ;
      RECT 8.32 1.12 11.105 1.135 ;
      RECT 9.2 1.135 11.105 1.29 ;
      RECT 9.2 1.29 10.085 1.45 ;
      RECT 10.835 1.29 11.105 1.8 ;
      RECT 2.055 2.31 5.775 2.46 ;
      RECT 3.155 2.46 5.775 2.48 ;
      RECT 5.215 1.47 5.385 2.31 ;
      RECT 5.605 2.48 5.775 2.89 ;
      RECT 5.215 1.3 5.785 1.47 ;
      RECT 5.605 2.89 6.445 3.06 ;
      RECT 5.535 0.595 5.785 1.3 ;
      RECT 1.375 2.905 2.225 3.075 ;
      RECT 2.055 2.46 2.225 2.905 ;
      RECT 2.055 2.29 3.545 2.31 ;
      RECT 3.155 2.48 3.545 2.96 ;
      RECT 3.375 0.81 3.545 2.29 ;
      RECT 3 0.35 3.545 0.81 ;
      RECT 1.375 2.46 1.545 2.905 ;
      RECT 0.085 2.29 1.545 2.46 ;
      RECT 0.085 2.46 0.445 2.98 ;
      RECT 0.085 0.42 0.6 0.75 ;
      RECT 0.085 0.75 0.255 2.29 ;
      RECT 4.165 1.81 4.965 2.14 ;
      RECT 4.555 1.01 4.725 1.81 ;
      RECT 4.065 0.84 4.725 1.01 ;
      RECT 4.065 0.35 4.395 0.84 ;
      RECT 6.65 2.72 6.98 2.98 ;
      RECT 6.55 2.55 6.98 2.72 ;
      RECT 6.55 1.91 6.72 2.55 ;
      RECT 6.55 1.74 8.26 1.91 ;
      RECT 7.93 1.91 8.26 1.955 ;
      RECT 6.55 1.685 6.72 1.74 ;
      RECT 7.93 1.645 8.26 1.74 ;
      RECT 6.295 1.515 6.72 1.685 ;
      RECT 6.295 0.595 6.465 1.515 ;
      RECT 13.265 1.32 13.975 1.65 ;
      RECT 12.155 0.255 13.435 0.425 ;
      RECT 13.265 0.425 13.435 1.32 ;
      RECT 12.45 2.12 12.7 2.845 ;
      RECT 11.615 1.805 12.7 2.12 ;
      RECT 11.615 1.725 12.485 1.805 ;
      RECT 12.155 0.425 12.485 1.725 ;
      RECT 2.875 0.98 3.205 1.99 ;
      RECT 0 -0.085 14.4 0.085 ;
      RECT 13.605 0.085 13.775 1.15 ;
      RECT 1.09 0.085 1.42 0.81 ;
      RECT 2.17 0.085 2.5 0.81 ;
      RECT 3.715 0.085 3.885 1.01 ;
      RECT 4.585 0.085 4.915 0.67 ;
      RECT 7.22 0.085 7.47 0.795 ;
      RECT 8.66 0.085 8.91 0.77 ;
      RECT 11.655 0.085 11.985 0.985 ;
      RECT 0 3.245 14.4 3.415 ;
      RECT 13.54 1.82 13.79 3.245 ;
      RECT 7.695 2.885 8.025 3.245 ;
      RECT 3.715 2.65 4.045 3.245 ;
      RECT 5.105 2.65 5.435 3.245 ;
      RECT 0.955 2.63 1.205 3.245 ;
      RECT 2.395 2.63 2.645 3.245 ;
      RECT 11.495 2.325 12.28 3.245 ;
      RECT 9.575 1.96 9.905 3.245 ;
  END
END scs8ls_edfxbp_1

MACRO scs8ls_edfxtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.075 1.55 12.405 2.98 ;
        RECT 12.075 1.13 12.345 1.55 ;
        RECT 12.015 0.35 12.345 1.13 ;
    END
    ANTENNADIFFAREA 0.5189 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.45 1.18 3.78 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.98 0.805 1.99 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END D

  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515 1.11 1.845 1.44 ;
    END
    ANTENNAGATEAREA 0.285 ;
  END DE

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12.96 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12.96 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 11.675 1.58 11.845 1.75 ;
      RECT 2.555 1.58 2.725 1.75 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
    LAYER met1 ;
      RECT 2.495 1.735 2.785 1.78 ;
      RECT 2.495 1.595 11.905 1.735 ;
      RECT 11.615 1.735 11.905 1.78 ;
      RECT 2.495 1.55 2.785 1.595 ;
      RECT 11.615 1.55 11.905 1.595 ;
    LAYER li1 ;
      RECT 3.1 2.12 3.475 2.31 ;
      RECT 3.1 2.31 5.61 2.48 ;
      RECT 3.1 2.48 3.475 2.62 ;
      RECT 5.44 2.48 5.61 2.52 ;
      RECT 5.13 1.65 5.3 2.31 ;
      RECT 5.44 2.52 6.245 2.69 ;
      RECT 5.13 1.48 5.655 1.65 ;
      RECT 5.995 2.69 6.245 2.98 ;
      RECT 5.325 0.595 5.655 1.48 ;
      RECT 1.365 2.905 2.215 3.075 ;
      RECT 1.365 2.35 1.535 2.905 ;
      RECT 2.045 2.12 2.215 2.905 ;
      RECT 0.085 2.18 1.535 2.35 ;
      RECT 2.045 1.95 3.27 2.12 ;
      RECT 3.1 0.875 3.27 1.95 ;
      RECT 2.79 0.415 3.27 0.875 ;
      RECT 0.085 2.35 0.435 2.98 ;
      RECT 0.085 0.34 0.53 0.81 ;
      RECT 0.085 0.81 0.255 2.18 ;
      RECT 6.945 2.41 9.8 2.58 ;
      RECT 6.945 2.33 7.115 2.41 ;
      RECT 9.63 1.725 9.8 2.41 ;
      RECT 6.755 2 7.115 2.33 ;
      RECT 9.63 1.545 10.065 1.725 ;
      RECT 5.825 2.14 6.245 2.3 ;
      RECT 5.47 1.97 6.245 2.14 ;
      RECT 5.47 1.82 5.995 1.97 ;
      RECT 5.825 0.425 5.995 1.82 ;
      RECT 4.765 0.255 6.96 0.425 ;
      RECT 4.765 0.425 5.095 1.13 ;
      RECT 6.79 0.425 6.96 0.935 ;
      RECT 6.505 0.935 7.76 1.105 ;
      RECT 6.505 1.105 6.96 1.31 ;
      RECT 7.59 0.425 7.76 0.935 ;
      RECT 7.59 0.255 8.44 0.425 ;
      RECT 8.27 0.425 8.44 0.935 ;
      RECT 8.27 0.935 9.28 1.105 ;
      RECT 9.11 1.105 9.28 1.205 ;
      RECT 9.11 1.205 10.605 1.375 ;
      RECT 9.11 1.375 9.46 1.55 ;
      RECT 10.275 1.375 10.605 1.585 ;
      RECT 0 -0.085 12.96 0.085 ;
      RECT 12.515 0.085 12.845 1.13 ;
      RECT 2 0.085 2.33 0.875 ;
      RECT 3.44 0.085 3.61 1.01 ;
      RECT 4.335 0.085 4.585 1.13 ;
      RECT 7.17 0.085 7.42 0.765 ;
      RECT 8.61 0.085 8.86 0.765 ;
      RECT 10.35 0.085 11.31 0.665 ;
      RECT 1.02 0.085 1.35 0.6 ;
      RECT 0 3.245 12.96 3.415 ;
      RECT 12.605 1.82 12.855 3.245 ;
      RECT 7.41 2.75 7.74 3.245 ;
      RECT 8.505 2.75 8.835 3.245 ;
      RECT 3.67 2.65 4 3.245 ;
      RECT 5.02 2.65 5.27 3.245 ;
      RECT 10.845 2.525 11.385 3.245 ;
      RECT 0.945 2.52 1.195 3.245 ;
      RECT 2.385 2.29 2.635 3.245 ;
      RECT 0.975 1.61 2.385 1.78 ;
      RECT 1.705 1.78 1.875 2.735 ;
      RECT 2.055 1.385 2.385 1.61 ;
      RECT 0.975 0.77 1.82 0.94 ;
      RECT 1.57 0.415 1.82 0.77 ;
      RECT 0.975 1.78 1.305 2.01 ;
      RECT 0.975 0.94 1.305 1.61 ;
      RECT 9.97 2.095 10.22 3 ;
      RECT 9.97 1.925 10.405 2.095 ;
      RECT 10.235 1.755 10.945 1.925 ;
      RECT 10.775 1.335 10.945 1.755 ;
      RECT 10.775 1.005 11.505 1.335 ;
      RECT 9.45 0.835 10.945 1.005 ;
      RECT 9.45 0.35 9.78 0.835 ;
      RECT 3.95 1.47 4.9 2.14 ;
      RECT 3.95 1.01 4.12 1.47 ;
      RECT 3.79 0.35 4.12 1.01 ;
      RECT 11.555 2.32 11.885 2.95 ;
      RECT 10.665 2.095 11.885 2.32 ;
      RECT 11.645 1.55 11.885 2.095 ;
      RECT 11.675 0.81 11.845 1.55 ;
      RECT 11.49 0.335 11.845 0.81 ;
      RECT 2.555 1.045 2.93 1.78 ;
      RECT 6.415 2.52 6.775 2.98 ;
      RECT 6.415 1.8 6.585 2.52 ;
      RECT 6.165 1.63 8.03 1.8 ;
      RECT 7.7 1.8 8.03 1.83 ;
      RECT 7.7 1.615 8.03 1.63 ;
      RECT 6.165 0.765 6.335 1.63 ;
      RECT 6.165 0.595 6.62 0.765 ;
      RECT 7.945 2.07 8.44 2.24 ;
      RECT 8.27 1.605 8.44 2.07 ;
      RECT 8.27 1.445 8.94 1.605 ;
      RECT 7.13 1.275 8.94 1.445 ;
      RECT 7.13 1.445 7.46 1.46 ;
      RECT 7.93 0.595 8.1 1.275 ;
  END
END scs8ls_edfxtp_1

MACRO scs8ls_einvn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455 1.43 1.315 1.76 ;
        RECT 1.085 1.76 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.327 ;
  END TEB

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.765 1.95 2.315 2.98 ;
        RECT 2.145 1.18 2.315 1.95 ;
        RECT 1.77 0.48 2.315 1.18 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END Z

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.35 1.975 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.39 2.1 0.72 2.58 ;
      RECT 0.11 1.93 0.72 2.1 ;
      RECT 0.11 0.56 0.77 1.25 ;
      RECT 0.11 0.255 0.78 0.56 ;
      RECT 0.11 1.25 0.28 1.93 ;
      RECT 0 3.245 2.4 3.415 ;
      RECT 0.925 1.95 1.255 3.245 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 0.95 0.085 1.28 1.26 ;
    LAYER mcon ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_einvn_1

MACRO scs8ls_einvn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.425 0.77 2.755 1.13 ;
        RECT 2.465 1.13 2.755 1.82 ;
        RECT 2.465 1.82 2.795 2.735 ;
    END
    ANTENNADIFFAREA 0.5469 ;
  END Z

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 0.81 3.255 1.55 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A

  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.12 0.55 2.13 ;
    END
    ANTENNAGATEAREA 0.495 ;
  END TEB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.015 2.905 3.245 3.075 ;
      RECT 2.965 1.82 3.245 2.905 ;
      RECT 1.115 1.99 1.4 2.98 ;
      RECT 1.115 1.82 2.295 1.99 ;
      RECT 2.015 1.99 2.295 2.905 ;
      RECT 2.075 0.35 3.2 0.6 ;
      RECT 1.135 0.98 2.245 1.15 ;
      RECT 2.075 0.6 2.245 0.98 ;
      RECT 1.135 0.35 1.385 0.98 ;
      RECT 0.56 2.3 0.89 2.98 ;
      RECT 0.72 1.65 0.89 2.3 ;
      RECT 0.72 1.32 1.16 1.65 ;
      RECT 0.72 0.81 0.89 1.32 ;
      RECT 0.56 0.35 0.89 0.81 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 0.13 0.085 0.38 0.81 ;
      RECT 1.565 0.085 1.895 0.79 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 0.11 2.3 0.36 3.245 ;
      RECT 1.58 2.16 1.815 3.245 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_einvn_2

MACRO scs8ls_einvn_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.55 3.815 1.72 ;
        RECT 3.485 1.72 4.715 1.89 ;
        RECT 3.615 1.13 3.815 1.55 ;
        RECT 3.485 1.89 3.815 2.735 ;
        RECT 4.385 1.89 4.715 2.735 ;
        RECT 3.615 1.01 3.865 1.13 ;
        RECT 3.615 0.77 4.655 1.01 ;
        RECT 4.485 0.595 4.655 0.77 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END Z

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.035 1.18 5.155 1.55 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A

  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.3 0.455 1.78 ;
    END
    ANTENNAGATEAREA 0.951 ;
  END TEB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.185 0.255 5.165 0.425 ;
      RECT 4.835 0.425 5.165 1.01 ;
      RECT 3.185 0.425 4.305 0.6 ;
      RECT 1.465 1.14 3.435 1.31 ;
      RECT 3.185 0.6 3.435 1.14 ;
      RECT 1.465 0.35 1.635 1.14 ;
      RECT 2.325 0.35 2.495 1.14 ;
      RECT 0.625 1.31 0.955 2.98 ;
      RECT 0.625 1.13 1.295 1.31 ;
      RECT 0.545 0.3 1.295 1.13 ;
      RECT 3.035 2.905 5.165 3.075 ;
      RECT 4.915 1.82 5.165 2.905 ;
      RECT 4.015 2.06 4.185 2.905 ;
      RECT 3.035 1.65 3.285 2.905 ;
      RECT 1.185 1.48 3.285 1.65 ;
      RECT 1.185 1.65 1.435 2.98 ;
      RECT 2.085 1.65 2.335 2.98 ;
      RECT 0 3.245 5.28 3.415 ;
      RECT 0.175 1.95 0.425 3.245 ;
      RECT 1.635 1.82 1.885 3.245 ;
      RECT 2.535 1.82 2.865 3.245 ;
      RECT 0 -0.085 5.28 0.085 ;
      RECT 0.115 0.085 0.365 1.13 ;
      RECT 1.815 0.085 2.145 0.97 ;
      RECT 2.675 0.085 3.005 0.97 ;
    LAYER mcon ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_einvn_4

MACRO scs8ls_einvn_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.55 5.725 1.78 ;
        RECT 5.555 1.78 5.725 1.95 ;
        RECT 5.455 1.13 5.725 1.55 ;
        RECT 5.555 1.95 8.555 2.12 ;
        RECT 5.455 1.01 8.505 1.13 ;
        RECT 5.555 2.12 5.725 2.735 ;
        RECT 6.425 2.12 6.755 2.735 ;
        RECT 7.325 2.12 7.655 2.735 ;
        RECT 8.225 2.12 8.555 2.735 ;
        RECT 6.315 1.13 8.505 1.18 ;
        RECT 5.455 0.77 6.645 1.01 ;
        RECT 7.325 0.615 7.495 1.01 ;
        RECT 8.175 0.615 8.505 1.01 ;
    END
    ANTENNADIFFAREA 2.3324 ;
  END Z

  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.435 1.63 ;
    END
    ANTENNAGATEAREA 1.623 ;
  END TEB

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.995 1.35 8.995 1.78 ;
    END
    ANTENNAGATEAREA 2.232 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 5.025 2.905 9.005 3.075 ;
      RECT 8.755 1.95 9.005 2.905 ;
      RECT 5.925 2.29 6.255 2.905 ;
      RECT 6.955 2.29 7.125 2.905 ;
      RECT 7.855 2.29 8.025 2.905 ;
      RECT 4.025 2.12 4.355 2.98 ;
      RECT 4.025 1.835 4.495 1.95 ;
      RECT 1.175 1.665 4.495 1.835 ;
      RECT 1.175 1.835 1.425 2.98 ;
      RECT 2.125 1.835 2.375 2.98 ;
      RECT 3.075 1.835 3.325 2.98 ;
      RECT 5.025 2.12 5.355 2.905 ;
      RECT 4.025 1.95 5.355 2.12 ;
      RECT 5.105 0.255 9.005 0.425 ;
      RECT 8.675 0.425 9.005 1.13 ;
      RECT 5.105 0.425 7.145 0.6 ;
      RECT 6.815 0.6 7.145 0.825 ;
      RECT 7.675 0.425 8.005 0.825 ;
      RECT 1.525 1.38 4.415 1.47 ;
      RECT 1.525 1.3 5.275 1.38 ;
      RECT 4.165 1.21 5.275 1.3 ;
      RECT 1.525 0.35 1.695 1.3 ;
      RECT 2.305 0.35 2.555 1.3 ;
      RECT 3.235 0.35 3.485 1.3 ;
      RECT 5.105 0.6 5.275 1.21 ;
      RECT 4.165 0.35 4.415 1.21 ;
      RECT 0.615 1.335 0.945 2.98 ;
      RECT 0.615 1.13 1.355 1.335 ;
      RECT 0.685 0.325 1.355 1.13 ;
      RECT 0 3.245 9.12 3.415 ;
      RECT 4.525 2.29 4.855 3.245 ;
      RECT 1.625 2.005 1.955 3.245 ;
      RECT 2.575 2.005 2.905 3.245 ;
      RECT 3.525 2.005 3.855 3.245 ;
      RECT 0.115 1.82 0.445 3.245 ;
      RECT 0 -0.085 9.12 0.085 ;
      RECT 0.175 0.085 0.505 0.99 ;
      RECT 1.875 0.085 2.125 1.13 ;
      RECT 2.735 0.085 3.065 1.13 ;
      RECT 3.665 0.085 3.995 1.13 ;
      RECT 4.595 0.085 4.925 1.04 ;
    LAYER mcon ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
  END
END scs8ls_einvn_8

MACRO scs8ls_einvp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945 1.3 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955 2.275 2.285 2.98 ;
        RECT 1.605 1.95 2.285 2.275 ;
        RECT 1.605 1.13 1.775 1.95 ;
        RECT 1.605 0.96 2.285 1.13 ;
        RECT 1.955 0.35 2.285 0.96 ;
    END
    ANTENNADIFFAREA 0.5059 ;
  END Z

  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.44 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END TE

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.105 2.745 0.89 3.075 ;
      RECT 0.105 2.01 0.88 2.745 ;
      RECT 0.105 0.41 0.94 1.06 ;
      RECT 0.105 1.06 0.275 2.01 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 1.135 0.085 1.42 1.13 ;
      RECT 0 3.245 2.4 3.415 ;
      RECT 1.085 2.02 1.415 3.245 ;
    LAYER mcon ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_einvp_1

MACRO scs8ls_einvp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.48 0.26 2.81 0.67 ;
    END
    ANTENNAGATEAREA 0.381 ;
  END TE

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.435 1.55 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.18 0.92 2.735 ;
        RECT 0.67 0.625 0.92 1.18 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END Z

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.415 1.14 2.745 2.98 ;
      RECT 2.415 0.84 2.8 1.14 ;
      RECT 1.1 1.14 2.21 1.31 ;
      RECT 1.1 0.425 1.27 1.14 ;
      RECT 1.95 0.35 2.21 1.14 ;
      RECT 0.16 0.255 1.27 0.425 ;
      RECT 0.16 0.425 0.49 1.01 ;
      RECT 0.115 2.905 1.265 3.075 ;
      RECT 1.095 1.65 1.265 2.905 ;
      RECT 1.095 1.48 2.165 1.65 ;
      RECT 1.915 1.65 2.165 2.98 ;
      RECT 0.115 1.82 0.365 2.905 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.915 2.3 3.245 3.245 ;
      RECT 1.465 1.82 1.715 3.245 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.98 0.085 3.245 1.01 ;
      RECT 1.45 0.085 1.78 0.97 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_einvp_2

MACRO scs8ls_einvp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.43 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 2.12 1.895 2.735 ;
        RECT 0.615 1.95 1.895 2.12 ;
        RECT 0.615 2.12 0.945 2.735 ;
        RECT 1.615 1.18 1.895 1.95 ;
        RECT 0.615 1.01 1.945 1.18 ;
        RECT 0.615 0.66 0.945 1.01 ;
        RECT 1.615 0.66 1.945 1.01 ;
    END
    ANTENNADIFFAREA 1.2219 ;
  END Z

  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405 1.18 5.65 1.3 ;
        RECT 4.98 1.3 5.65 1.63 ;
    END
    ANTENNAGATEAREA 0.723 ;
  END TE

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.115 2.905 2.395 3.075 ;
      RECT 2.065 1.81 2.395 2.905 ;
      RECT 2.065 1.64 4.175 1.81 ;
      RECT 3.015 1.81 3.265 2.98 ;
      RECT 3.925 1.81 4.175 2.98 ;
      RECT 0.115 1.95 0.445 2.905 ;
      RECT 1.115 2.29 1.365 2.905 ;
      RECT 2.115 1.3 4.445 1.47 ;
      RECT 2.115 0.425 2.445 1.3 ;
      RECT 3.115 0.35 3.445 1.3 ;
      RECT 4.115 0.35 4.445 1.3 ;
      RECT 0.115 0.255 2.445 0.425 ;
      RECT 0.115 0.425 0.445 1.13 ;
      RECT 1.115 0.425 1.445 0.8 ;
      RECT 4.395 1.82 5.195 2.98 ;
      RECT 4.615 0.35 5.005 1.13 ;
      RECT 4.395 2.98 4.785 2.99 ;
      RECT 4.395 1.64 4.785 1.82 ;
      RECT 4.615 1.13 4.785 1.64 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 2.565 1.98 2.815 3.245 ;
      RECT 3.465 1.98 3.725 3.245 ;
      RECT 5.395 1.82 5.645 3.245 ;
      RECT 2.615 0.085 2.945 1.13 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 3.615 0.085 3.945 1.13 ;
      RECT 5.175 0.085 5.505 1.01 ;
    LAYER mcon ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_einvp_4

MACRO scs8ls_einvp_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.41 1.18 3.46 1.55 ;
    END
    ANTENNAGATEAREA 2.232 ;
  END A

  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.435 1.18 8.995 1.41 ;
        RECT 8.435 1.41 8.765 1.55 ;
    END
    ANTENNAGATEAREA 1.167 ;
  END TE

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.705 1.55 4.195 1.72 ;
        RECT 0.56 1.72 4.195 1.89 ;
        RECT 3.705 1.01 3.875 1.55 ;
        RECT 0.56 1.89 0.89 2.735 ;
        RECT 1.46 1.89 1.79 2.735 ;
        RECT 2.36 1.89 2.69 2.735 ;
        RECT 3.26 1.89 3.59 2.735 ;
        RECT 0.625 0.84 3.875 1.01 ;
        RECT 0.625 0.615 0.875 0.84 ;
        RECT 1.545 0.615 1.875 0.84 ;
        RECT 2.545 0.615 2.875 0.84 ;
        RECT 3.545 0.595 3.875 0.84 ;
    END
    ANTENNADIFFAREA 2.3282 ;
  END Z

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.11 2.905 3.96 3.075 ;
      RECT 3.79 2.23 3.96 2.905 ;
      RECT 3.79 2.06 4.94 2.23 ;
      RECT 4.69 2.23 4.94 2.98 ;
      RECT 4.69 1.72 4.94 2.06 ;
      RECT 4.69 1.55 7.56 1.72 ;
      RECT 5.51 1.72 5.76 2.98 ;
      RECT 6.41 1.72 6.66 2.98 ;
      RECT 7.31 1.72 7.56 2.98 ;
      RECT 0.11 1.82 0.375 2.905 ;
      RECT 1.07 2.06 1.275 2.905 ;
      RECT 1.97 2.06 2.19 2.905 ;
      RECT 2.875 2.06 3.075 2.905 ;
      RECT 8.235 2.965 8.565 2.98 ;
      RECT 7.775 1.82 8.565 2.965 ;
      RECT 8.055 0.35 8.505 1.01 ;
      RECT 7.775 1.615 8.225 1.82 ;
      RECT 8.055 1.01 8.225 1.615 ;
      RECT 4.055 1.21 7.885 1.38 ;
      RECT 4.055 0.425 4.225 1.21 ;
      RECT 4.905 0.35 5.155 1.21 ;
      RECT 5.845 0.35 6.015 1.21 ;
      RECT 6.705 0.35 6.955 1.21 ;
      RECT 7.635 0.35 7.885 1.21 ;
      RECT 0.115 0.255 4.225 0.425 ;
      RECT 0.115 0.425 0.445 1.01 ;
      RECT 1.045 0.425 1.375 0.67 ;
      RECT 2.045 0.425 2.375 0.67 ;
      RECT 3.045 0.425 3.375 0.67 ;
      RECT 0 3.245 9.12 3.415 ;
      RECT 4.16 2.4 4.49 3.245 ;
      RECT 5.14 1.89 5.31 3.245 ;
      RECT 5.96 1.89 6.21 3.245 ;
      RECT 6.86 1.89 7.11 3.245 ;
      RECT 8.765 1.82 9.015 3.245 ;
      RECT 4.405 0.085 4.735 1.04 ;
      RECT 0 -0.085 9.12 0.085 ;
      RECT 5.335 0.085 5.665 1.04 ;
      RECT 6.195 0.085 6.525 1.04 ;
      RECT 7.125 0.085 7.455 1.04 ;
      RECT 8.675 0.085 8.935 1.01 ;
    LAYER mcon ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
  END
END scs8ls_einvp_8

MACRO scs8ls_fa_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.35 0.365 1.13 ;
        RECT 0.085 1.13 0.255 1.82 ;
        RECT 0.085 1.82 0.355 2.98 ;
    END
    ANTENNADIFFAREA 0.5301 ;
  END SUM

  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.21 0.35 8.54 1.13 ;
        RECT 8.285 1.13 8.54 2.98 ;
    END
    ANTENNADIFFAREA 0.519 ;
  END COUT

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.8 1.32 7.47 1.78 ;
    END
    ANTENNAGATEAREA 0.984 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.38 1.105 4.71 1.455 ;
        RECT 4.38 1.09 5.98 1.105 ;
        RECT 5.81 1.105 5.98 1.32 ;
        RECT 1.045 0.935 5.98 1.09 ;
        RECT 5.81 1.32 6.21 1.575 ;
        RECT 1.045 1.09 1.215 1.22 ;
        RECT 3.3 1.09 3.63 1.455 ;
        RECT 1.045 0.92 4.71 0.935 ;
        RECT 0.885 1.22 1.215 1.54 ;
    END
    ANTENNAGATEAREA 0.984 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.535 1.595 5.185 1.735 ;
        RECT 1.535 1.735 1.825 1.78 ;
        RECT 3.935 1.735 4.225 1.78 ;
        RECT 4.895 1.735 5.185 1.78 ;
        RECT 1.535 1.55 1.825 1.595 ;
        RECT 3.935 1.55 4.225 1.595 ;
        RECT 4.895 1.55 5.185 1.595 ;
    END
    ANTENNAGATEAREA 0.738 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.604 LAYER met1 ;
  END CIN

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 5.665 2.255 5.95 2.755 ;
      RECT 5.665 2.085 7.32 2.255 ;
      RECT 7 2.255 7.32 2.83 ;
      RECT 6.99 1.95 7.32 2.085 ;
      RECT 4.925 1.575 5.155 1.78 ;
      RECT 4.925 1.275 5.64 1.575 ;
      RECT 3.84 1.26 4.195 1.78 ;
      RECT 2.61 2.46 2.86 2.755 ;
      RECT 2.61 2.29 3.93 2.46 ;
      RECT 3.6 2.46 3.93 2.755 ;
      RECT 2.61 1.965 2.86 2.29 ;
      RECT 2.48 0.58 3.91 0.75 ;
      RECT 2.48 0.42 2.89 0.58 ;
      RECT 3.58 0.42 3.91 0.58 ;
      RECT 2.08 2.12 2.41 2.755 ;
      RECT 1.055 1.95 2.41 2.12 ;
      RECT 1.055 1.88 1.225 1.95 ;
      RECT 2.08 1.745 2.41 1.95 ;
      RECT 0.535 1.71 1.225 1.88 ;
      RECT 0.535 0.58 2.27 0.75 ;
      RECT 1.94 0.355 2.27 0.58 ;
      RECT 0.535 1.63 0.705 1.71 ;
      RECT 0.425 1.3 0.705 1.63 ;
      RECT 0.535 0.75 0.705 1.3 ;
      RECT 1.565 1.575 1.795 1.78 ;
      RECT 1.565 1.26 2.115 1.575 ;
      RECT 0 -0.085 8.64 0.085 ;
      RECT 0.625 0.085 0.98 0.41 ;
      RECT 3.07 0.085 3.4 0.41 ;
      RECT 4.08 0.085 4.555 0.71 ;
      RECT 6.83 0.085 7.08 0.47 ;
      RECT 7.78 0.085 8.03 0.77 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 3.08 2.63 3.41 3.245 ;
      RECT 6.12 2.5 6.825 3.245 ;
      RECT 4.105 2.305 4.435 3.245 ;
      RECT 0.555 2.05 0.885 3.245 ;
      RECT 7.755 1.82 8.085 3.245 ;
      RECT 6.15 0.98 8.04 1.15 ;
      RECT 7.71 1.15 8.04 1.55 ;
      RECT 5.325 1.745 6.55 1.915 ;
      RECT 6.38 1.15 6.55 1.745 ;
      RECT 6.15 0.765 6.32 0.98 ;
      RECT 5.045 0.595 6.32 0.765 ;
      RECT 3.03 1.795 3.2 1.95 ;
      RECT 2.58 1.625 3.2 1.795 ;
      RECT 2.58 1.575 2.75 1.625 ;
      RECT 2.325 1.26 2.75 1.575 ;
      RECT 5.07 2.12 5.495 2.755 ;
      RECT 3.03 1.95 5.495 2.12 ;
      RECT 5.325 1.915 5.495 1.95 ;
      RECT 5.045 0.435 5.375 0.595 ;
      RECT 6.49 0.64 7.59 0.81 ;
      RECT 7.26 0.48 7.59 0.64 ;
      RECT 6.49 0.425 6.66 0.64 ;
      RECT 5.555 0.255 6.66 0.425 ;
    LAYER mcon ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 1.58 5.125 1.75 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 1.58 4.165 1.75 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 1.58 1.765 1.75 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_fa_1

MACRO scs8ls_fa_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.22 1.82 8.575 2.98 ;
        RECT 8.405 1.15 8.575 1.82 ;
        RECT 8.245 0.375 8.575 1.15 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END SUM

  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.985 1.82 7.555 2.15 ;
        RECT 7.385 1.085 7.555 1.82 ;
        RECT 7.105 0.915 7.555 1.085 ;
    END
    ANTENNADIFFAREA 0.6496 ;
  END COUT

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.92 0.835 2.15 ;
        RECT 0.665 1.575 0.835 1.92 ;
        RECT 0.665 1.245 1.165 1.575 ;
    END
    ANTENNAGATEAREA 1.044 ;
  END B

  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.055 1.95 4.535 2.105 ;
        RECT 2.055 2.105 4.195 2.12 ;
        RECT 3.375 1.935 4.535 1.95 ;
        RECT 2.055 1.575 2.225 1.95 ;
        RECT 3.375 2.12 4.195 2.15 ;
        RECT 4.365 1.915 4.535 1.935 ;
        RECT 3.375 1.575 3.545 1.935 ;
        RECT 1.715 1.26 2.225 1.575 ;
        RECT 4.365 1.745 5.635 1.915 ;
        RECT 3.215 1.26 3.545 1.575 ;
        RECT 5.305 1.26 5.635 1.745 ;
    END
    ANTENNAGATEAREA 0.783 ;
  END CIN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
    END
  END vpwr

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.095 1.595 6.625 1.735 ;
        RECT 0.095 1.735 0.385 1.78 ;
        RECT 0.095 1.55 0.385 1.595 ;
        RECT 2.495 1.735 2.785 1.78 ;
        RECT 3.935 1.735 4.225 1.78 ;
        RECT 6.335 1.735 6.625 1.78 ;
        RECT 2.495 1.55 2.785 1.595 ;
        RECT 3.935 1.55 4.225 1.595 ;
        RECT 6.335 1.55 6.625 1.595 ;
    END
    ANTENNAGATEAREA 1.044 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.683 LAYER met1 ;
  END A

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.965 1.26 4.525 1.575 ;
      RECT 3.965 1.575 4.195 1.765 ;
      RECT 2.525 1.575 2.755 1.78 ;
      RECT 2.525 1.26 3.005 1.575 ;
      RECT 0.115 1.075 0.445 1.13 ;
      RECT 0.115 0.905 1.205 1.075 ;
      RECT 1.035 0.75 1.205 0.905 ;
      RECT 0.115 0.375 0.445 0.905 ;
      RECT 1.035 0.42 1.81 0.75 ;
      RECT 3.48 0.58 4.97 0.75 ;
      RECT 4.5 0.42 4.97 0.58 ;
      RECT 3.48 0.375 3.81 0.58 ;
      RECT 0.095 2.32 1.545 2.49 ;
      RECT 1.215 2.49 1.545 2.755 ;
      RECT 1.215 2.085 1.545 2.32 ;
      RECT 0.095 2.49 0.445 2.91 ;
      RECT 0.095 1.95 0.425 2.32 ;
      RECT 6.765 1.255 7.165 1.585 ;
      RECT 1.375 0.92 6.935 1.09 ;
      RECT 6.765 1.09 6.935 1.255 ;
      RECT 1.375 1.09 1.545 1.745 ;
      RECT 1.715 1.915 1.885 2.29 ;
      RECT 1.375 1.745 1.885 1.915 ;
      RECT 1.715 2.29 2.185 2.62 ;
      RECT 1.98 0.375 2.31 0.92 ;
      RECT 4.765 1.09 5.095 1.575 ;
      RECT 3.405 2.49 3.735 2.755 ;
      RECT 3.405 2.32 4.825 2.49 ;
      RECT 4.495 2.49 4.825 2.755 ;
      RECT 4.495 2.275 4.825 2.32 ;
      RECT 7.88 1.32 8.235 1.65 ;
      RECT 5.005 2.32 8.05 2.49 ;
      RECT 7.88 1.65 8.05 2.32 ;
      RECT 7.88 0.745 8.05 1.32 ;
      RECT 5.14 0.575 8.05 0.745 ;
      RECT 5.005 2.49 5.335 2.755 ;
      RECT 5.005 2.085 5.335 2.32 ;
      RECT 5.14 0.745 5.47 0.75 ;
      RECT 5.14 0.375 5.47 0.575 ;
      RECT 6.265 1.35 6.595 1.78 ;
      RECT 0.105 1.3 0.435 1.78 ;
      RECT 0 3.245 9.12 3.415 ;
      RECT 8.75 1.82 9 3.245 ;
      RECT 7.53 2.73 8.05 3.245 ;
      RECT 6.535 2.66 6.865 3.245 ;
      RECT 0.615 2.66 1.01 3.245 ;
      RECT 2.825 2.29 3.155 3.245 ;
      RECT 3.905 2.66 4.29 3.245 ;
      RECT 0 -0.085 9.12 0.085 ;
      RECT 8.755 0.085 9.005 1.155 ;
      RECT 7.615 0.085 8.065 0.405 ;
      RECT 0.615 0.085 0.865 0.735 ;
      RECT 2.8 0.085 3.31 0.705 ;
      RECT 3.99 0.085 4.32 0.41 ;
      RECT 6.47 0.085 6.925 0.405 ;
    LAYER mcon ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 1.58 0.325 1.75 ;
      RECT 3.995 1.58 4.165 1.75 ;
      RECT 2.555 1.58 2.725 1.75 ;
      RECT 6.395 1.58 6.565 1.75 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
  END
END scs8ls_fa_2

MACRO scs8ls_fa_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 11.04 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.245 0.835 1.78 ;
    END
    ANTENNAGATEAREA 1.044 ;
  END A

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.195 2.01 8.525 2.98 ;
        RECT 7.245 1.84 8.525 2.01 ;
        RECT 7.245 2.01 7.575 2.98 ;
        RECT 8.285 1.17 8.525 1.84 ;
        RECT 7.265 0.92 8.615 1.17 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END SUM

  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.165 1.55 10.435 1.82 ;
        RECT 9.145 1.82 10.435 1.99 ;
        RECT 10.165 1.15 10.425 1.55 ;
        RECT 9.145 1.99 9.475 2.98 ;
        RECT 10.095 1.99 10.435 2.98 ;
        RECT 9.305 0.98 10.425 1.15 ;
        RECT 9.305 0.39 9.555 0.98 ;
        RECT 10.165 0.39 10.425 0.98 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END COUT

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.915 1.55 6.595 1.72 ;
        RECT 4.45 1.72 6.595 1.745 ;
        RECT 5.915 1.26 6.34 1.55 ;
        RECT 2.48 1.745 6.595 1.78 ;
        RECT 2.48 1.78 6.085 1.89 ;
        RECT 3.95 1.26 4.28 1.745 ;
        RECT 2.48 1.245 2.81 1.745 ;
        RECT 2.48 1.89 4.62 1.915 ;
        RECT 2.48 1.915 2.65 1.95 ;
        RECT 1.665 1.95 2.65 2.12 ;
        RECT 1.665 1.575 1.835 1.95 ;
        RECT 1.345 1.26 1.835 1.575 ;
    END
    ANTENNAGATEAREA 1.044 ;
  END B

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.04 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.04 3.575 ;
    END
  END vpwr

  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2.015 1.225 5.665 1.365 ;
        RECT 2.015 1.365 2.305 1.41 ;
        RECT 2.015 1.18 2.305 1.225 ;
        RECT 2.975 1.365 3.265 1.41 ;
        RECT 5.375 1.365 5.665 1.41 ;
        RECT 2.975 1.18 3.265 1.225 ;
        RECT 5.375 1.18 5.665 1.225 ;
    END
    ANTENNAGATEAREA 0.783 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.604 LAYER met1 ;
  END CIN

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.005 1.26 3.74 1.575 ;
      RECT 3.005 1.18 3.215 1.26 ;
      RECT 0.985 2.63 2.005 2.96 ;
      RECT 0.985 2.255 1.155 2.63 ;
      RECT 0.115 2.085 1.155 2.255 ;
      RECT 0.115 2.255 0.445 2.98 ;
      RECT 0.115 1.95 0.445 2.085 ;
      RECT 0.115 0.75 0.445 1.075 ;
      RECT 0.115 0.67 1.495 0.75 ;
      RECT 0.115 0.58 1.965 0.67 ;
      RECT 0.115 0.35 0.445 0.58 ;
      RECT 1.325 0.35 1.965 0.58 ;
      RECT 3.725 0.58 4.915 0.75 ;
      RECT 3.725 0.35 3.975 0.58 ;
      RECT 4.665 0.35 4.915 0.58 ;
      RECT 8.965 1.32 9.955 1.65 ;
      RECT 6.255 0.58 9.135 0.75 ;
      RECT 8.965 0.75 9.135 1.32 ;
      RECT 5.085 0.255 6.425 0.425 ;
      RECT 6.255 0.425 6.425 0.58 ;
      RECT 1.005 1.09 1.175 1.745 ;
      RECT 1.325 1.915 1.495 2.29 ;
      RECT 1.005 1.745 1.495 1.915 ;
      RECT 1.005 1.01 1.835 1.09 ;
      RECT 2.135 0.35 2.465 0.84 ;
      RECT 2.21 2.46 2.54 2.755 ;
      RECT 1.325 2.29 2.54 2.46 ;
      RECT 1.665 0.84 3.555 0.92 ;
      RECT 1.005 0.92 5.255 1.01 ;
      RECT 3.385 1.01 5.255 1.09 ;
      RECT 5.085 0.425 5.255 0.92 ;
      RECT 4.93 1.09 5.255 1.22 ;
      RECT 4.93 1.22 5.26 1.55 ;
      RECT 3.67 2.255 4 2.755 ;
      RECT 3.67 2.085 5.07 2.255 ;
      RECT 4.74 2.255 5.07 2.755 ;
      RECT 6.905 1.34 8.105 1.67 ;
      RECT 5.24 2.12 6.425 2.23 ;
      RECT 5.24 2.06 7.075 2.12 ;
      RECT 6.255 1.95 7.075 2.06 ;
      RECT 6.905 1.67 7.075 1.95 ;
      RECT 6.905 1.09 7.075 1.34 ;
      RECT 5.915 1.01 7.075 1.09 ;
      RECT 5.425 0.92 7.075 1.01 ;
      RECT 5.425 0.84 6.085 0.92 ;
      RECT 5.24 2.23 5.57 2.755 ;
      RECT 5.425 0.595 5.675 0.84 ;
      RECT 5.43 1.18 5.745 1.55 ;
      RECT 2.005 1.18 2.275 1.78 ;
      RECT 0 3.245 11.04 3.415 ;
      RECT 10.625 1.82 10.875 3.245 ;
      RECT 8.725 1.82 8.975 3.245 ;
      RECT 4.17 2.425 4.57 3.245 ;
      RECT 6.795 2.29 7.045 3.245 ;
      RECT 3.17 2.085 3.5 3.245 ;
      RECT 7.775 2.18 8.025 3.245 ;
      RECT 9.675 2.16 9.925 3.245 ;
      RECT 0.645 2.425 0.815 3.245 ;
      RECT 0 -0.085 11.04 0.085 ;
      RECT 10.595 0.085 10.925 1.17 ;
      RECT 7.775 0.085 8.105 0.41 ;
      RECT 8.795 0.085 9.125 0.41 ;
      RECT 0.625 0.085 1.155 0.41 ;
      RECT 3.175 0.085 3.505 0.67 ;
      RECT 4.155 0.085 4.485 0.41 ;
      RECT 6.755 0.085 7.085 0.41 ;
      RECT 9.735 0.085 9.985 0.81 ;
    LAYER mcon ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 1.21 3.205 1.38 ;
      RECT 5.435 1.21 5.605 1.38 ;
      RECT 2.075 1.21 2.245 1.38 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
  END
END scs8ls_fa_4

MACRO scs8ls_fah_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 13.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.145 1.18 9.475 1.55 ;
    END
    ANTENNAGATEAREA 0.723 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.072 LAYER li1 ;
  END B

  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505 0.4 2.075 0.73 ;
        RECT 0.665 0.73 1.675 0.9 ;
        RECT 0.665 0.9 0.835 1.95 ;
        RECT 0.665 1.95 1.155 2.12 ;
        RECT 0.985 2.12 1.155 2.905 ;
        RECT 0.985 2.905 2.645 3.075 ;
        RECT 2.315 2.875 2.645 2.905 ;
    END
    ANTENNADIFFAREA 0.67485 ;
    ANTENNAPARTIALMETALSIDEAREA 1.117 LAYER li1 ;
  END COUT

  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 0.54 0.445 2.98 ;
    END
    ANTENNADIFFAREA 0.5376 ;
    ANTENNAPARTIALMETALSIDEAREA 0.215 LAYER li1 ;
  END SUM

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.41 1.335 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.072 LAYER li1 ;
  END CI

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.82 1.47 13.49 1.8 ;
    END
    ANTENNAGATEAREA 0.492 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.132 LAYER li1 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.92 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 11.91 0.79 12.805 0.96 ;
      RECT 12.475 0.35 12.805 0.79 ;
      RECT 9.28 1.805 10.475 2.395 ;
      RECT 9.645 0.96 9.975 1.805 ;
      RECT 3.495 2.025 4 2.115 ;
      RECT 3.005 1.855 4 2.025 ;
      RECT 3.005 1.58 3.445 1.855 ;
      RECT 3.275 1.185 3.445 1.58 ;
      RECT 3.275 0.935 3.605 1.185 ;
      RECT 5.405 1.705 5.635 2.15 ;
      RECT 5.405 1.375 5.885 1.705 ;
      RECT 6.845 1.55 7.075 1.78 ;
      RECT 6.845 1.38 7.065 1.55 ;
      RECT 6.735 0.71 7.065 1.38 ;
      RECT 8.17 2.905 11.74 3.075 ;
      RECT 11.385 1.13 11.74 2.905 ;
      RECT 11.405 0.35 11.74 1.13 ;
      RECT 8.17 1.88 8.61 2.905 ;
      RECT 8.17 1.21 8.34 1.88 ;
      RECT 8.17 0.96 8.635 1.21 ;
      RECT 6.33 2.49 6.66 2.64 ;
      RECT 5.045 2.32 6.66 2.49 ;
      RECT 6.33 2.29 6.66 2.32 ;
      RECT 5.045 1.425 5.215 2.32 ;
      RECT 4.88 1.265 5.215 1.425 ;
      RECT 3.775 1.095 5.215 1.265 ;
      RECT 3.775 0.765 3.945 1.095 ;
      RECT 2.935 0.595 3.945 0.765 ;
      RECT 2.935 0.765 3.105 1.24 ;
      RECT 2.5 1.24 3.105 1.41 ;
      RECT 2.5 1.41 2.83 1.635 ;
      RECT 4.205 2.455 4.535 2.735 ;
      RECT 3.155 2.365 4.535 2.455 ;
      RECT 1.845 2.285 4.535 2.365 ;
      RECT 1.845 2.195 3.325 2.285 ;
      RECT 4.205 2.1 4.535 2.285 ;
      RECT 1.845 1.07 2.175 2.195 ;
      RECT 1.845 0.9 2.765 1.07 ;
      RECT 2.595 0.425 2.765 0.9 ;
      RECT 2.595 0.255 4.285 0.425 ;
      RECT 4.115 0.425 4.285 0.755 ;
      RECT 4.115 0.755 6.215 0.765 ;
      RECT 4.115 0.765 5.045 0.925 ;
      RECT 5.885 0.765 6.215 0.865 ;
      RECT 4.875 0.595 6.215 0.755 ;
      RECT 6.395 1.55 6.595 1.78 ;
      RECT 6.395 0.67 6.565 1.55 ;
      RECT 3.46 2.905 7 3.075 ;
      RECT 3.46 2.795 3.63 2.905 ;
      RECT 4.705 2.73 6.125 2.905 ;
      RECT 6.83 2.12 7 2.905 ;
      RECT 2.815 2.705 3.63 2.795 ;
      RECT 4.705 1.765 4.875 2.73 ;
      RECT 6.055 1.95 7 2.12 ;
      RECT 1.325 2.625 3.63 2.705 ;
      RECT 4.17 1.685 4.875 1.765 ;
      RECT 6.055 1.205 6.225 1.95 ;
      RECT 1.325 2.535 2.985 2.625 ;
      RECT 3.67 1.595 4.875 1.685 ;
      RECT 5.385 1.035 6.225 1.205 ;
      RECT 3.67 1.435 4.34 1.595 ;
      RECT 5.385 0.935 5.715 1.035 ;
      RECT 1.325 2.705 1.675 2.735 ;
      RECT 1.325 1.95 1.675 2.535 ;
      RECT 1.505 1.24 1.675 1.95 ;
      RECT 1.13 1.07 1.675 1.24 ;
      RECT 7.235 0.62 10.315 0.79 ;
      RECT 10.145 0.79 10.315 1.22 ;
      RECT 10.145 1.22 10.475 1.55 ;
      RECT 7.17 1.95 7.5 2.925 ;
      RECT 7.33 1.13 7.5 1.95 ;
      RECT 7.235 0.79 7.565 1.13 ;
      RECT 8.805 0.79 8.975 1.38 ;
      RECT 7.235 0.425 7.565 0.62 ;
      RECT 8.51 1.38 8.975 1.71 ;
      RECT 4.455 0.255 7.565 0.425 ;
      RECT 4.455 0.425 4.705 0.585 ;
      RECT 13.47 1.97 13.83 2.98 ;
      RECT 13.66 1.3 13.83 1.97 ;
      RECT 12.25 1.13 13.83 1.3 ;
      RECT 13.475 0.35 13.83 1.13 ;
      RECT 12.25 1.3 12.58 1.55 ;
      RECT 10.985 1.78 11.155 2.735 ;
      RECT 10.985 1.55 11.215 1.78 ;
      RECT 10.985 0.425 11.155 1.55 ;
      RECT 8.895 0.255 11.155 0.425 ;
      RECT 8.895 0.425 9.385 0.45 ;
      RECT 8.78 2.565 10.815 2.735 ;
      RECT 10.645 1.05 10.815 2.565 ;
      RECT 10.485 0.595 10.815 1.05 ;
      RECT 8.78 1.88 9.11 2.565 ;
      RECT 0 3.245 13.92 3.415 ;
      RECT 13.05 1.97 13.3 3.245 ;
      RECT 2.935 2.965 3.29 3.245 ;
      RECT 11.95 2.33 12.29 3.245 ;
      RECT 7.67 1.765 8 3.245 ;
      RECT 11.95 2.11 12.22 2.33 ;
      RECT 0.645 2.29 0.815 3.245 ;
      RECT 0 -0.085 13.92 0.085 ;
      RECT 2.255 0.085 2.425 0.73 ;
      RECT 7.745 0.085 8.075 0.45 ;
      RECT 11.915 0.085 12.245 0.62 ;
      RECT 12.975 0.085 13.305 0.96 ;
      RECT 0.62 0.085 0.95 0.56 ;
      RECT 12.52 2.16 12.85 2.98 ;
      RECT 12.39 1.97 12.85 2.16 ;
      RECT 12.39 1.94 12.65 1.97 ;
      RECT 11.91 1.72 12.65 1.94 ;
      RECT 11.91 0.96 12.08 1.72 ;
    LAYER mcon ;
      RECT 10.245 1.95 10.415 2.12 ;
      RECT 9.885 1.95 10.055 2.12 ;
      RECT 8.84 1.95 9.01 2.12 ;
      RECT 6.395 1.58 6.565 1.75 ;
      RECT 3.035 1.58 3.205 1.75 ;
      RECT 11.015 1.58 11.185 1.75 ;
      RECT 6.875 1.58 7.045 1.75 ;
      RECT 5.435 1.95 5.605 2.12 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 12.435 1.95 12.605 2.12 ;
    LAYER met1 ;
      RECT 2.975 1.735 3.265 1.78 ;
      RECT 2.975 1.595 6.625 1.735 ;
      RECT 6.335 1.735 6.625 1.78 ;
      RECT 2.975 1.55 3.265 1.595 ;
      RECT 6.335 1.55 6.625 1.595 ;
      RECT 9.825 2.105 10.475 2.15 ;
      RECT 9.825 1.965 12.665 2.105 ;
      RECT 12.375 2.105 12.665 2.15 ;
      RECT 9.825 1.92 10.475 1.965 ;
      RECT 12.375 1.92 12.665 1.965 ;
      RECT 6.815 1.735 7.105 1.78 ;
      RECT 6.815 1.595 11.245 1.735 ;
      RECT 10.955 1.735 11.245 1.78 ;
      RECT 6.815 1.55 7.105 1.595 ;
      RECT 10.955 1.55 11.245 1.595 ;
      RECT 5.375 2.105 5.665 2.15 ;
      RECT 5.375 1.965 9.07 2.105 ;
      RECT 8.78 2.105 9.07 2.15 ;
      RECT 5.375 1.92 5.665 1.965 ;
      RECT 8.78 1.92 9.07 1.965 ;
  END
END scs8ls_fah_1

MACRO scs8ls_dfstp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 11.04 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.315 1.18 1.795 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475 0.98 0.805 1.99 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.5 0.35 10.935 1.05 ;
        RECT 10.685 1.05 10.935 2.98 ;
    END
    ANTENNADIFFAREA 0.5301 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.04 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.04 3.575 ;
    END
  END vpwr

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.375 1.965 8.545 2.105 ;
        RECT 8.255 2.105 8.545 2.15 ;
        RECT 8.255 1.92 8.545 1.965 ;
        RECT 5.375 2.105 5.665 2.15 ;
        RECT 5.375 1.92 5.665 1.965 ;
    END
    ANTENNAGATEAREA 0.252 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.205 LAYER met1 ;
  END SETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 5.435 1.95 5.605 2.12 ;
      RECT 8.315 1.95 8.485 2.12 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
    LAYER li1 ;
      RECT 8.185 1.13 8.515 2.14 ;
      RECT 0 3.245 11.04 3.415 ;
      RECT 5.535 2.66 5.785 3.245 ;
      RECT 7.77 2.65 7.94 3.245 ;
      RECT 8.665 2.65 8.915 3.245 ;
      RECT 0.555 2.57 0.885 3.245 ;
      RECT 1.54 2.57 1.87 3.245 ;
      RECT 3.95 2.425 4.23 3.245 ;
      RECT 10.155 1.82 10.485 3.245 ;
      RECT 0 -0.085 11.04 0.085 ;
      RECT 0.545 0.085 0.795 0.81 ;
      RECT 1.615 0.085 1.785 1.01 ;
      RECT 4.065 0.085 4.455 0.68 ;
      RECT 5.62 0.085 5.95 1.03 ;
      RECT 7.87 0.085 8.76 0.6 ;
      RECT 10 0.085 10.33 1.03 ;
      RECT 3.08 2.295 3.415 2.735 ;
      RECT 3.245 1.02 3.415 2.295 ;
      RECT 3.245 0.85 4.095 1.02 ;
      RECT 3.925 1.02 4.095 1.345 ;
      RECT 3.245 0.415 3.575 0.85 ;
      RECT 3.925 1.345 6.065 1.515 ;
      RECT 4.805 1.515 6.065 1.545 ;
      RECT 4.805 1.215 6.065 1.345 ;
      RECT 2.83 1.435 3.075 2.105 ;
      RECT 2.905 0.425 3.075 1.435 ;
      RECT 1.965 0.255 3.075 0.425 ;
      RECT 1.965 0.425 2.295 1.09 ;
      RECT 4.74 2.32 5.025 2.735 ;
      RECT 4.74 1.915 4.91 2.32 ;
      RECT 4.055 1.745 4.91 1.915 ;
      RECT 4.055 1.685 4.385 1.745 ;
      RECT 2.07 2.905 3.755 3.075 ;
      RECT 2.07 2.4 2.32 2.905 ;
      RECT 3.585 2.255 3.755 2.905 ;
      RECT 3.585 2.085 4.57 2.255 ;
      RECT 4.4 2.255 4.57 2.905 ;
      RECT 3.585 1.435 3.755 2.085 ;
      RECT 4.4 2.905 5.365 3.075 ;
      RECT 5.195 2.49 5.365 2.905 ;
      RECT 5.195 2.32 5.975 2.49 ;
      RECT 5.805 1.885 5.975 2.32 ;
      RECT 5.805 1.715 6.405 1.885 ;
      RECT 6.235 1.45 6.405 1.715 ;
      RECT 6.235 1.12 6.645 1.45 ;
      RECT 6.235 0.425 6.405 1.12 ;
      RECT 6.235 0.255 7.325 0.425 ;
      RECT 7.155 0.425 7.325 1.97 ;
      RECT 6.98 1.97 7.325 2.14 ;
      RECT 6.98 2.14 7.26 2.355 ;
      RECT 4.265 1.03 4.625 1.175 ;
      RECT 4.265 0.86 5.01 1.03 ;
      RECT 4.625 0.57 5.01 0.86 ;
      RECT 5.08 1.82 5.635 2.15 ;
      RECT 9.635 1.22 10.515 1.55 ;
      RECT 9.635 1.55 9.965 2.875 ;
      RECT 9.635 0.86 9.82 1.22 ;
      RECT 9.49 0.35 9.82 0.86 ;
      RECT 6.475 2.625 7.6 2.98 ;
      RECT 7.43 2.48 7.6 2.625 ;
      RECT 6.475 2.05 6.81 2.625 ;
      RECT 7.43 2.31 9.105 2.48 ;
      RECT 6.575 1.8 6.81 2.05 ;
      RECT 8.14 2.48 8.47 2.93 ;
      RECT 8.775 1.37 9.105 2.31 ;
      RECT 6.575 1.63 6.985 1.8 ;
      RECT 6.815 0.925 6.985 1.63 ;
      RECT 6.575 0.595 6.985 0.925 ;
      RECT 9.115 2.65 9.445 2.98 ;
      RECT 9.275 1.2 9.445 2.65 ;
      RECT 9.09 1.03 9.445 1.2 ;
      RECT 9.09 0.96 9.26 1.03 ;
      RECT 7.495 0.79 9.26 0.96 ;
      RECT 7.495 0.96 7.73 1.555 ;
      RECT 8.93 0.35 9.26 0.79 ;
      RECT 0.105 2.23 1.76 2.4 ;
      RECT 1.59 2.06 2.66 2.23 ;
      RECT 2.49 2.23 2.66 2.295 ;
      RECT 2.485 0.925 2.66 2.06 ;
      RECT 2.49 2.295 2.91 2.735 ;
      RECT 2.485 0.595 2.735 0.925 ;
      RECT 0.105 2.4 0.355 2.98 ;
      RECT 0.105 0.81 0.275 2.23 ;
      RECT 0.105 0.35 0.365 0.81 ;
      RECT 0.975 1.89 1.42 2.06 ;
      RECT 0.975 1.72 2.315 1.89 ;
      RECT 1.985 1.26 2.315 1.72 ;
      RECT 0.975 0.35 1.435 1.01 ;
      RECT 0.975 1.01 1.145 1.72 ;
  END
END scs8ls_dfstp_1

MACRO scs8ls_dfstp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.685 1.82 11.465 2.15 ;
        RECT 11.155 2.15 11.465 2.98 ;
        RECT 11.295 1.13 11.465 1.82 ;
        RECT 11.1 0.35 11.465 1.13 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475 0.98 0.805 1.99 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.315 1.18 1.775 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12 3.575 ;
    END
  END vpwr

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.855 1.965 8.545 2.105 ;
        RECT 8.255 2.105 8.545 2.15 ;
        RECT 8.255 1.92 8.545 1.965 ;
        RECT 5.855 2.105 6.145 2.15 ;
        RECT 5.855 1.92 6.145 1.965 ;
    END
    ANTENNAGATEAREA 0.252 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.869 LAYER met1 ;
  END SETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.915 1.95 6.085 2.12 ;
      RECT 8.315 1.95 8.485 2.12 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
    LAYER li1 ;
      RECT 0 3.245 12 3.415 ;
      RECT 11.635 1.82 11.885 3.245 ;
      RECT 4.07 2.91 4.24 3.245 ;
      RECT 8.1 2.72 8.43 3.245 ;
      RECT 5.86 2.66 6.11 3.245 ;
      RECT 9.11 2.66 9.44 3.245 ;
      RECT 0.565 2.53 0.895 3.245 ;
      RECT 1.575 2.53 1.905 3.245 ;
      RECT 4.07 2.58 4.575 2.91 ;
      RECT 10.655 2.32 10.985 3.245 ;
      RECT 4.425 1.05 4.77 1.23 ;
      RECT 4.425 0.88 5.16 1.05 ;
      RECT 4.77 0.57 5.16 0.88 ;
      RECT 2.785 1.38 3.115 2.05 ;
      RECT 2.945 0.425 3.115 1.38 ;
      RECT 2.045 0.255 3.115 0.425 ;
      RECT 2.045 0.425 2.215 1.13 ;
      RECT 5.085 2.32 5.35 2.72 ;
      RECT 5.085 2.07 5.255 2.32 ;
      RECT 4.23 1.74 5.255 2.07 ;
      RECT 7.83 1.24 8.145 2.13 ;
      RECT 7.83 1.07 9.89 1.24 ;
      RECT 9.64 1.24 9.89 2.98 ;
      RECT 9.53 0.635 9.89 1.07 ;
      RECT 2.105 2.89 3.795 3.06 ;
      RECT 3.625 2.41 3.795 2.89 ;
      RECT 2.105 2.4 2.275 2.89 ;
      RECT 3.625 2.24 4.915 2.41 ;
      RECT 4.745 2.41 4.915 2.89 ;
      RECT 3.625 1.38 3.915 2.24 ;
      RECT 4.745 2.89 5.69 3.06 ;
      RECT 5.52 2.49 5.69 2.89 ;
      RECT 5.52 2.32 6.585 2.49 ;
      RECT 6.415 1.45 6.585 2.32 ;
      RECT 6.415 1.12 6.96 1.45 ;
      RECT 6.415 0.45 6.585 1.12 ;
      RECT 6.415 0.28 7.66 0.45 ;
      RECT 7.49 0.45 7.66 1.98 ;
      RECT 7.29 1.98 7.66 2.15 ;
      RECT 7.29 2.15 7.59 2.38 ;
      RECT 0.975 1.89 1.455 2.02 ;
      RECT 0.975 1.72 2.275 1.89 ;
      RECT 1.945 1.3 2.275 1.72 ;
      RECT 0.975 0.35 1.435 1.01 ;
      RECT 0.975 1.01 1.145 1.72 ;
      RECT 3.115 2.26 3.455 2.72 ;
      RECT 3.285 1.21 3.455 2.26 ;
      RECT 3.285 1.04 4.255 1.21 ;
      RECT 4.085 1.21 4.255 1.4 ;
      RECT 3.285 0.4 3.615 1.04 ;
      RECT 4.085 1.4 6.245 1.57 ;
      RECT 4.95 1.22 6.245 1.4 ;
      RECT 5.915 1.215 6.245 1.22 ;
      RECT 6.82 2.73 7.47 2.98 ;
      RECT 6.82 2.55 7.93 2.73 ;
      RECT 7.76 2.49 8.88 2.55 ;
      RECT 6.82 1.79 7.07 2.55 ;
      RECT 8.63 2.55 8.88 2.98 ;
      RECT 7.76 2.32 9.47 2.49 ;
      RECT 6.82 1.62 7.32 1.79 ;
      RECT 9.14 1.615 9.47 2.32 ;
      RECT 7.15 0.95 7.32 1.62 ;
      RECT 6.825 0.62 7.32 0.95 ;
      RECT 10.09 1.3 11.125 1.63 ;
      RECT 10.09 1.63 10.45 2.86 ;
      RECT 10.09 0.45 10.42 1.3 ;
      RECT 5.425 1.79 6.115 2.15 ;
      RECT 0.115 2.23 1.795 2.36 ;
      RECT 0.115 2.19 2.615 2.23 ;
      RECT 2.445 2.23 2.615 2.26 ;
      RECT 1.625 2.06 2.615 2.19 ;
      RECT 2.445 2.26 2.945 2.72 ;
      RECT 2.445 0.925 2.615 2.06 ;
      RECT 2.445 0.595 2.775 0.925 ;
      RECT 0.115 2.36 0.365 2.98 ;
      RECT 0.115 0.765 0.285 2.19 ;
      RECT 0.115 0.395 0.365 0.765 ;
      RECT 8.315 1.48 8.73 2.15 ;
      RECT 0 -0.085 12 0.085 ;
      RECT 11.635 0.085 11.885 1.13 ;
      RECT 0.545 0.085 0.795 0.765 ;
      RECT 1.615 0.085 1.865 1.01 ;
      RECT 4.27 0.085 4.6 0.71 ;
      RECT 5.65 0.085 6.245 1.03 ;
      RECT 8.525 0.085 9.36 0.9 ;
      RECT 10.6 0.085 10.93 1.13 ;
  END
END scs8ls_dfstp_2

MACRO scs8ls_dfstp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.605 1.15 12.835 1.82 ;
        RECT 11.175 1.82 12.835 2.08 ;
        RECT 10.68 0.98 12.835 1.15 ;
        RECT 12.125 2.08 12.835 2.15 ;
        RECT 11.175 2.08 11.455 2.98 ;
        RECT 10.68 0.35 11.01 0.98 ;
        RECT 12.015 0.35 12.345 0.98 ;
        RECT 12.125 2.15 12.355 2.98 ;
    END
    ANTENNADIFFAREA 1.1197 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475 0.98 0.805 1.99 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.315 1.18 1.775 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12.96 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12.96 3.575 ;
    END
  END vpwr

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.375 1.595 8.545 1.735 ;
        RECT 8.255 1.735 8.545 1.78 ;
        RECT 8.255 1.55 8.545 1.595 ;
        RECT 5.375 1.735 5.665 1.78 ;
        RECT 5.375 1.55 5.665 1.595 ;
    END
    ANTENNAGATEAREA 0.252 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.205 LAYER met1 ;
  END SETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 1.58 5.605 1.75 ;
      RECT 8.315 1.58 8.485 1.75 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
    LAYER li1 ;
      RECT 0.115 2.24 1.795 2.41 ;
      RECT 1.625 2.07 2.615 2.24 ;
      RECT 2.445 2.24 2.615 2.295 ;
      RECT 2.445 0.925 2.615 2.07 ;
      RECT 2.445 2.295 2.945 2.735 ;
      RECT 2.445 0.595 2.775 0.925 ;
      RECT 0.115 2.41 0.365 2.96 ;
      RECT 0.115 0.81 0.285 2.24 ;
      RECT 0.115 0.35 0.365 0.81 ;
      RECT 8.185 1.18 8.515 1.85 ;
      RECT 0 -0.085 12.96 0.085 ;
      RECT 12.515 0.085 12.845 0.81 ;
      RECT 0.545 0.085 0.795 0.81 ;
      RECT 1.615 0.085 1.865 1.01 ;
      RECT 4.025 0.085 4.42 0.6 ;
      RECT 5.67 0.085 6 1.03 ;
      RECT 7.935 0.085 8.95 0.67 ;
      RECT 10.18 0.085 10.51 1.13 ;
      RECT 11.18 0.085 11.845 0.8 ;
      RECT 0 3.245 12.96 3.415 ;
      RECT 12.525 2.32 12.855 3.245 ;
      RECT 3.985 2.755 4.155 3.245 ;
      RECT 7.885 2.65 8.055 3.245 ;
      RECT 8.78 2.65 9.03 3.245 ;
      RECT 0.565 2.58 0.895 3.245 ;
      RECT 1.575 2.58 1.905 3.245 ;
      RECT 5.68 2.435 5.94 3.245 ;
      RECT 9.755 1.82 10.005 3.245 ;
      RECT 10.725 1.82 11.005 3.245 ;
      RECT 3.985 2.505 4.345 2.755 ;
      RECT 11.625 2.25 11.955 3.245 ;
      RECT 4.305 0.95 4.59 1.23 ;
      RECT 4.305 0.78 5.05 0.95 ;
      RECT 4.59 0.62 5.05 0.78 ;
      RECT 2.785 1.455 3.115 2.125 ;
      RECT 2.945 0.425 3.115 1.455 ;
      RECT 2.045 0.255 3.115 0.425 ;
      RECT 2.045 0.425 2.215 1.13 ;
      RECT 4.855 2.295 5.17 2.735 ;
      RECT 4.855 1.995 5.025 2.295 ;
      RECT 4.115 1.74 5.025 1.995 ;
      RECT 2.105 2.905 3.795 3.075 ;
      RECT 2.105 2.41 2.275 2.905 ;
      RECT 3.625 2.335 3.795 2.905 ;
      RECT 3.625 2.165 4.685 2.335 ;
      RECT 4.515 2.335 4.685 2.905 ;
      RECT 3.625 1.47 3.795 2.165 ;
      RECT 4.515 2.905 5.51 3.075 ;
      RECT 5.34 2.265 5.51 2.905 ;
      RECT 5.34 2.095 6.475 2.265 ;
      RECT 6.305 1.45 6.475 2.095 ;
      RECT 6.305 1.12 6.695 1.45 ;
      RECT 6.305 0.425 6.475 1.12 ;
      RECT 6.305 0.255 7.375 0.425 ;
      RECT 7.205 0.425 7.375 2.02 ;
      RECT 7.045 2.02 7.375 2.31 ;
      RECT 10.205 1.49 11.995 1.65 ;
      RECT 9.68 1.32 11.995 1.49 ;
      RECT 10.205 1.65 10.535 2.7 ;
      RECT 9.68 0.35 10.01 1.32 ;
      RECT 0.975 1.89 1.455 2.07 ;
      RECT 0.975 1.72 2.275 1.89 ;
      RECT 1.945 1.35 2.275 1.72 ;
      RECT 0.975 0.34 1.435 1.01 ;
      RECT 0.975 1.01 1.145 1.72 ;
      RECT 3.115 2.295 3.455 2.735 ;
      RECT 3.285 1.3 3.455 2.295 ;
      RECT 3.285 1.13 4.135 1.3 ;
      RECT 3.965 1.3 4.135 1.4 ;
      RECT 3.285 0.35 3.535 1.13 ;
      RECT 3.965 1.4 5.025 1.57 ;
      RECT 4.77 1.37 5.025 1.4 ;
      RECT 4.77 1.2 6.135 1.37 ;
      RECT 5.805 1.37 6.135 1.49 ;
      RECT 4.77 1.12 5.025 1.2 ;
      RECT 6.59 2.65 7.265 2.98 ;
      RECT 6.67 2.48 7.715 2.65 ;
      RECT 7.545 2.31 9.11 2.48 ;
      RECT 6.67 1.79 6.84 2.48 ;
      RECT 8.255 2.48 8.585 2.98 ;
      RECT 8.78 1.37 9.11 2.31 ;
      RECT 6.67 1.62 7.035 1.79 ;
      RECT 6.865 0.925 7.035 1.62 ;
      RECT 6.645 0.595 7.035 0.925 ;
      RECT 9.23 2.65 9.56 2.98 ;
      RECT 9.28 1.01 9.45 2.65 ;
      RECT 7.545 0.84 9.45 1.01 ;
      RECT 7.545 1.01 7.875 1.655 ;
      RECT 9.12 0.42 9.45 0.84 ;
      RECT 5.195 1.55 5.635 1.925 ;
  END
END scs8ls_dfstp_4

MACRO scs8ls_dfxbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.16 1.82 9.515 2.98 ;
        RECT 9.345 1.13 9.515 1.82 ;
        RECT 9.14 0.35 9.515 1.13 ;
    END
    ANTENNADIFFAREA 0.5357 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.665 2.03 8.07 2.98 ;
        RECT 7.9 1.13 8.07 2.03 ;
        RECT 7.64 0.35 8.07 1.13 ;
    END
    ANTENNADIFFAREA 0.5301 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.5 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.91 1.125 2.27 1.78 ;
        RECT 1.91 1.78 2.08 2.025 ;
        RECT 1.7 2.025 2.08 2.355 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 4.64 2.025 4.81 2.615 ;
      RECT 4.45 1.855 4.81 2.025 ;
      RECT 4.45 1.37 4.62 1.855 ;
      RECT 3.825 1.185 4.62 1.37 ;
      RECT 3.825 1.015 4.9 1.185 ;
      RECT 4.57 0.92 4.9 1.015 ;
      RECT 2.25 2.045 2.61 2.375 ;
      RECT 2.44 1.24 2.61 2.045 ;
      RECT 2.44 1.07 2.885 1.24 ;
      RECT 2.715 0.595 2.885 1.07 ;
      RECT 5.32 2.115 5.57 2.735 ;
      RECT 5.32 1.38 5.49 2.115 ;
      RECT 5.32 1.21 7.13 1.38 ;
      RECT 6.8 1.38 7.13 1.52 ;
      RECT 6.8 1.19 7.13 1.21 ;
      RECT 5.32 1.12 5.59 1.21 ;
      RECT 5.125 0.79 5.59 1.12 ;
      RECT 6.23 1.69 7.73 1.86 ;
      RECT 7.3 1.35 7.73 1.69 ;
      RECT 6.71 2.22 7.04 2.86 ;
      RECT 6.23 1.86 7.04 2.22 ;
      RECT 6.23 1.55 6.56 1.69 ;
      RECT 7.3 1.02 7.47 1.35 ;
      RECT 6.64 0.85 7.47 1.02 ;
      RECT 6.64 0.44 6.97 0.85 ;
      RECT 8.28 1.3 9.175 1.63 ;
      RECT 8.28 1.63 8.455 2.7 ;
      RECT 8.28 0.625 8.53 1.3 ;
      RECT 0.115 0.73 2.545 0.9 ;
      RECT 2.375 0.425 2.545 0.73 ;
      RECT 2.375 0.255 3.655 0.425 ;
      RECT 3.485 0.425 3.655 0.58 ;
      RECT 3.485 0.58 5.715 0.62 ;
      RECT 3.485 0.62 4.65 0.75 ;
      RECT 4.48 0.29 5.715 0.58 ;
      RECT 3.485 0.75 3.655 1.75 ;
      RECT 3.12 1.75 3.655 2.075 ;
      RECT 0.11 1.89 0.36 2.98 ;
      RECT 0.11 1.72 0.84 1.89 ;
      RECT 0.67 1.55 0.84 1.72 ;
      RECT 0.67 0.9 1.09 1.55 ;
      RECT 0.115 0.9 0.445 1.01 ;
      RECT 0.115 0.35 0.445 0.73 ;
      RECT 2.78 2.415 2.95 2.545 ;
      RECT 2.78 2.245 4.28 2.415 ;
      RECT 4.02 1.63 4.28 2.245 ;
      RECT 2.78 1.58 2.95 2.245 ;
      RECT 2.78 1.41 3.315 1.58 ;
      RECT 3.065 0.595 3.315 1.41 ;
      RECT 4.3 2.905 5.99 3.075 ;
      RECT 4.3 2.8 5.15 2.905 ;
      RECT 5.82 1.945 5.99 2.905 ;
      RECT 4.3 2.755 4.47 2.8 ;
      RECT 4.98 1.685 5.15 2.8 ;
      RECT 5.66 1.615 5.99 1.945 ;
      RECT 2.055 2.715 4.47 2.755 ;
      RECT 4.79 1.355 5.15 1.685 ;
      RECT 2.055 2.755 3.29 2.885 ;
      RECT 3.12 2.585 4.47 2.715 ;
      RECT 1.01 2.545 2.225 2.715 ;
      RECT 1.01 2.715 1.34 2.98 ;
      RECT 1.01 1.815 1.435 2.545 ;
      RECT 1.265 1.07 1.595 1.485 ;
      RECT 1.265 1.485 1.74 1.815 ;
      RECT 0 3.245 9.6 3.415 ;
      RECT 8.655 1.82 8.985 3.245 ;
      RECT 3.74 2.925 4.13 3.245 ;
      RECT 6.165 2.39 6.495 3.245 ;
      RECT 7.24 2.03 7.49 3.245 ;
      RECT 0.56 2.06 0.81 3.245 ;
      RECT 1.555 2.885 1.885 3.245 ;
      RECT 0 -0.085 9.6 0.085 ;
      RECT 8.71 0.085 8.96 1.13 ;
      RECT 1.855 0.085 2.205 0.56 ;
      RECT 3.98 0.085 4.31 0.41 ;
      RECT 6.08 0.085 6.41 1.04 ;
      RECT 7.14 0.085 7.47 0.68 ;
      RECT 0.625 0.085 1.005 0.56 ;
    LAYER mcon ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
  END
END scs8ls_dfxbp_1

MACRO scs8ls_dfxbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 11.04 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.14 1.82 10.505 2.98 ;
        RECT 10.335 1.13 10.505 1.82 ;
        RECT 10.165 0.35 10.505 1.13 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END QN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 1.125 2.375 1.78 ;
        RECT 1.985 1.78 2.155 2.025 ;
        RECT 1.825 2.025 2.155 2.355 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.145 1.55 8.515 2.07 ;
        RECT 8.145 0.37 8.45 1.55 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.585 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.04 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.04 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 5.375 1.79 5.705 2.625 ;
      RECT 5.375 1.67 7.585 1.79 ;
      RECT 6.375 1.79 7.585 1.96 ;
      RECT 5.375 1.62 6.545 1.67 ;
      RECT 6.015 0.95 6.185 1.62 ;
      RECT 5.785 0.7 6.185 0.95 ;
      RECT 7.16 2.24 9.015 2.41 ;
      RECT 8.685 1.32 9.015 2.24 ;
      RECT 7.16 2.41 7.49 2.98 ;
      RECT 7.16 2.13 7.925 2.24 ;
      RECT 7.755 1.5 7.925 2.13 ;
      RECT 6.715 1.33 7.925 1.5 ;
      RECT 6.715 1.17 7.465 1.33 ;
      RECT 7.215 0.37 7.465 1.17 ;
      RECT 0.115 0.73 2.53 0.9 ;
      RECT 2.36 0.425 2.53 0.73 ;
      RECT 2.36 0.255 3.64 0.425 ;
      RECT 3.47 0.425 3.64 0.78 ;
      RECT 3.47 0.78 4.815 0.95 ;
      RECT 3.47 0.95 3.64 1.75 ;
      RECT 4.645 0.53 4.815 0.78 ;
      RECT 3.225 1.75 3.64 2.065 ;
      RECT 4.645 0.255 6.24 0.53 ;
      RECT 5.445 0.53 5.615 1.17 ;
      RECT 5.445 1.17 5.845 1.45 ;
      RECT 0.115 1.89 0.445 2.98 ;
      RECT 0.115 1.72 0.925 1.89 ;
      RECT 0.755 1.55 0.925 1.72 ;
      RECT 0.755 1.01 1.1 1.55 ;
      RECT 0.115 0.9 1.1 1.01 ;
      RECT 0.115 0.35 0.445 0.73 ;
      RECT 4.535 2.18 4.865 2.455 ;
      RECT 4.645 1.45 4.815 2.18 ;
      RECT 3.81 1.12 4.815 1.45 ;
      RECT 2.885 2.285 4.325 2.455 ;
      RECT 4.155 1.96 4.325 2.285 ;
      RECT 2.885 1.58 3.055 2.285 ;
      RECT 4.155 1.63 4.475 1.96 ;
      RECT 2.885 1.41 3.3 1.58 ;
      RECT 3.05 0.595 3.3 1.41 ;
      RECT 2.325 2.205 2.715 2.455 ;
      RECT 2.545 1.24 2.715 2.205 ;
      RECT 2.545 1.07 2.87 1.24 ;
      RECT 2.7 0.595 2.87 1.07 ;
      RECT 1.095 2.625 5.205 2.795 ;
      RECT 5.035 2.795 6.205 2.965 ;
      RECT 5.035 1.45 5.205 2.625 ;
      RECT 5.875 1.96 6.205 2.795 ;
      RECT 4.985 1.12 5.275 1.45 ;
      RECT 1.095 2.795 1.345 2.98 ;
      RECT 1.095 1.815 1.44 2.625 ;
      RECT 1.27 1.485 1.815 1.815 ;
      RECT 1.27 1.07 1.6 1.485 ;
      RECT 9.235 1.3 10.165 1.63 ;
      RECT 9.235 1.63 9.485 2.86 ;
      RECT 9.235 0.54 9.51 1.3 ;
      RECT 0 -0.085 11.04 0.085 ;
      RECT 10.675 0.085 10.925 1.13 ;
      RECT 8.62 0.085 8.95 1.15 ;
      RECT 9.735 0.085 9.985 1.13 ;
      RECT 1.86 0.085 2.19 0.56 ;
      RECT 4.03 0.085 4.37 0.61 ;
      RECT 6.655 0.085 6.985 1 ;
      RECT 7.645 0.085 7.975 1.15 ;
      RECT 0.625 0.085 1.01 0.56 ;
      RECT 0 3.245 11.04 3.415 ;
      RECT 10.675 1.82 10.925 3.245 ;
      RECT 8.595 2.58 8.925 3.245 ;
      RECT 9.69 1.82 9.94 3.245 ;
      RECT 1.575 2.965 2.035 3.245 ;
      RECT 4 2.965 4.33 3.245 ;
      RECT 7.695 2.58 8.025 3.245 ;
      RECT 6.6 2.375 6.93 3.245 ;
      RECT 0.645 2.06 0.895 3.245 ;
    LAYER mcon ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
  END
END scs8ls_dfxbp_2

MACRO scs8ls_dfxtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.87 2.025 2.25 2.355 ;
        RECT 1.97 1.125 2.25 2.025 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.715 0.35 8.075 1.13 ;
        RECT 7.905 1.13 8.075 2.03 ;
        RECT 7.715 2.03 8.075 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.3 0.505 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 4.335 2.125 4.61 2.455 ;
      RECT 4.44 1.2 4.61 2.125 ;
      RECT 3.93 1.03 5 1.2 ;
      RECT 3.93 1.2 4.26 1.415 ;
      RECT 4.83 0.595 5 1.03 ;
      RECT 2.76 2.455 3.12 2.625 ;
      RECT 2.76 2.285 4.14 2.455 ;
      RECT 3.97 1.955 4.14 2.285 ;
      RECT 2.76 1.58 2.93 2.285 ;
      RECT 3.97 1.625 4.27 1.955 ;
      RECT 2.76 1.41 3.42 1.58 ;
      RECT 3.155 0.615 3.42 1.41 ;
      RECT 2.42 1.24 2.59 2.625 ;
      RECT 2.42 1.07 2.975 1.24 ;
      RECT 6.05 1.69 7.735 1.86 ;
      RECT 7.375 1.35 7.735 1.69 ;
      RECT 6.05 1.86 6.38 2.24 ;
      RECT 6.76 1.86 7.01 2.7 ;
      RECT 6.05 1.57 6.38 1.69 ;
      RECT 7.375 1.02 7.545 1.35 ;
      RECT 6.79 0.85 7.545 1.02 ;
      RECT 6.79 0.35 7.04 0.85 ;
      RECT 1.645 0.73 2.655 0.9 ;
      RECT 2.485 0.445 2.655 0.73 ;
      RECT 2.485 0.275 3.76 0.445 ;
      RECT 3.59 0.445 3.76 0.69 ;
      RECT 3.59 0.69 4.66 0.86 ;
      RECT 3.59 0.86 3.76 1.75 ;
      RECT 4.49 0.425 4.66 0.69 ;
      RECT 3.1 1.75 3.76 2.08 ;
      RECT 4.49 0.255 5.895 0.425 ;
      RECT 5.565 0.425 5.895 0.51 ;
      RECT 0.115 2.12 0.445 2.98 ;
      RECT 0.115 1.95 0.845 2.12 ;
      RECT 0.675 1.55 0.845 1.95 ;
      RECT 0.675 1.13 1.135 1.55 ;
      RECT 0.115 0.96 1.135 1.13 ;
      RECT 0.965 0.425 1.135 0.96 ;
      RECT 0.115 0.35 0.365 0.96 ;
      RECT 0.965 0.255 1.815 0.425 ;
      RECT 1.645 0.425 1.815 0.73 ;
      RECT 5.12 1.88 5.29 2.735 ;
      RECT 5.12 1.71 5.82 1.88 ;
      RECT 5.65 1.4 5.82 1.71 ;
      RECT 5.65 1.23 7.205 1.4 ;
      RECT 6.875 1.4 7.205 1.52 ;
      RECT 6.875 1.19 7.205 1.23 ;
      RECT 5.65 0.98 5.82 1.23 ;
      RECT 5.22 0.73 5.82 0.98 ;
      RECT 1.015 2.625 2.25 2.795 ;
      RECT 2.08 2.795 3.46 2.965 ;
      RECT 3.29 2.625 4.95 2.795 ;
      RECT 4.78 2.795 4.95 2.905 ;
      RECT 4.78 1.54 4.95 2.625 ;
      RECT 4.78 2.905 5.84 3.075 ;
      RECT 4.78 1.37 5.48 1.54 ;
      RECT 5.51 2.05 5.84 2.905 ;
      RECT 5.17 1.15 5.48 1.37 ;
      RECT 1.015 2.795 1.345 2.98 ;
      RECT 1.015 1.82 1.475 2.625 ;
      RECT 1.305 1.68 1.475 1.82 ;
      RECT 1.305 1.35 1.76 1.68 ;
      RECT 1.305 0.595 1.475 1.35 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 1.575 2.965 1.91 3.245 ;
      RECT 3.8 2.965 4.13 3.245 ;
      RECT 6.2 2.52 6.53 3.245 ;
      RECT 7.21 2.03 7.54 3.245 ;
      RECT 0.645 2.29 0.815 3.245 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 0.545 0.085 0.795 0.79 ;
      RECT 1.985 0.085 2.315 0.56 ;
      RECT 4.07 0.085 4.32 0.52 ;
      RECT 6.23 0.085 6.56 1.06 ;
      RECT 7.22 0.085 7.535 0.68 ;
    LAYER mcon ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
  END
END scs8ls_dfxtp_1

MACRO scs8ls_dfxtp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885 1.15 2.275 1.48 ;
        RECT 1.885 1.48 2.055 2.05 ;
        RECT 1.725 2.05 2.055 2.38 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.3 0.505 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.745 2.03 8.105 2.98 ;
        RECT 7.935 1.13 8.105 2.03 ;
        RECT 7.765 0.35 8.105 1.13 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 4.305 2.125 4.65 2.455 ;
      RECT 4.48 1.415 4.65 2.125 ;
      RECT 3.925 1.2 4.65 1.415 ;
      RECT 3.925 1.03 4.915 1.2 ;
      RECT 4.745 0.945 4.915 1.03 ;
      RECT 4.745 0.595 5.075 0.945 ;
      RECT 5.16 1.88 5.33 2.735 ;
      RECT 5.16 1.71 5.755 1.88 ;
      RECT 5.585 1.4 5.755 1.71 ;
      RECT 5.585 1.23 7.24 1.4 ;
      RECT 6.91 1.4 7.24 1.52 ;
      RECT 6.91 1.19 7.24 1.23 ;
      RECT 5.585 0.945 5.755 1.23 ;
      RECT 5.245 0.695 5.755 0.945 ;
      RECT 2.755 2.425 2.955 2.585 ;
      RECT 2.755 2.255 4.135 2.425 ;
      RECT 2.755 2.125 2.955 2.255 ;
      RECT 3.965 1.955 4.135 2.255 ;
      RECT 2.785 1.66 2.955 2.125 ;
      RECT 3.965 1.625 4.31 1.955 ;
      RECT 2.785 1.49 3.2 1.66 ;
      RECT 3.03 0.945 3.2 1.49 ;
      RECT 3.03 0.615 3.415 0.945 ;
      RECT 2.225 1.82 2.555 2.455 ;
      RECT 2.225 1.65 2.615 1.82 ;
      RECT 2.445 1.32 2.615 1.65 ;
      RECT 2.445 1.15 2.86 1.32 ;
      RECT 2.69 0.595 2.86 1.15 ;
      RECT 1.015 2.755 4.99 2.795 ;
      RECT 2.105 2.795 3.54 2.925 ;
      RECT 4.82 2.795 4.99 2.905 ;
      RECT 1.015 2.625 2.275 2.755 ;
      RECT 3.37 2.625 4.99 2.755 ;
      RECT 4.82 2.905 5.875 3.075 ;
      RECT 4.82 1.54 4.99 2.625 ;
      RECT 5.545 2.05 5.875 2.905 ;
      RECT 4.82 1.37 5.415 1.54 ;
      RECT 5.085 1.15 5.415 1.37 ;
      RECT 1.015 2.795 1.345 2.98 ;
      RECT 1.015 1.72 1.475 2.625 ;
      RECT 1.305 1.35 1.715 1.72 ;
      RECT 1.305 0.595 1.475 1.35 ;
      RECT 6.085 1.69 7.765 1.86 ;
      RECT 7.425 1.35 7.765 1.69 ;
      RECT 6.085 1.86 6.415 2.24 ;
      RECT 6.79 1.86 7.04 2.86 ;
      RECT 6.085 1.57 6.415 1.69 ;
      RECT 7.425 1.02 7.595 1.35 ;
      RECT 6.785 0.85 7.595 1.02 ;
      RECT 6.785 0.35 7.115 0.85 ;
      RECT 1.645 0.81 2.52 0.98 ;
      RECT 2.35 0.425 2.52 0.81 ;
      RECT 2.35 0.255 3.755 0.425 ;
      RECT 3.585 0.425 3.755 0.69 ;
      RECT 3.585 0.69 4.575 0.86 ;
      RECT 3.585 0.86 3.755 1.285 ;
      RECT 4.405 0.425 4.575 0.69 ;
      RECT 3.37 1.285 3.755 1.455 ;
      RECT 4.405 0.255 5.89 0.425 ;
      RECT 3.37 1.455 3.54 1.83 ;
      RECT 5.56 0.425 5.89 0.51 ;
      RECT 3.14 1.83 3.54 2.085 ;
      RECT 0.115 2.12 0.445 2.98 ;
      RECT 0.115 1.95 0.845 2.12 ;
      RECT 0.675 1.55 0.845 1.95 ;
      RECT 0.675 1.13 1.135 1.55 ;
      RECT 0.115 0.96 1.135 1.13 ;
      RECT 0.965 0.425 1.135 0.96 ;
      RECT 0.115 0.35 0.365 0.96 ;
      RECT 0.965 0.255 1.815 0.425 ;
      RECT 1.645 0.425 1.815 0.81 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 8.275 1.82 8.525 3.245 ;
      RECT 1.575 2.965 1.935 3.245 ;
      RECT 3.71 2.965 4.1 3.245 ;
      RECT 6.235 2.52 6.565 3.245 ;
      RECT 7.24 2.03 7.57 3.245 ;
      RECT 0.645 2.29 0.815 3.245 ;
      RECT 0 -0.085 8.64 0.085 ;
      RECT 8.275 0.085 8.525 1.13 ;
      RECT 0.545 0.085 0.795 0.79 ;
      RECT 1.985 0.085 2.18 0.64 ;
      RECT 3.985 0.085 4.235 0.52 ;
      RECT 6.225 0.085 6.555 1.06 ;
      RECT 7.3 0.085 7.595 0.68 ;
    LAYER mcon ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_dfxtp_2

MACRO scs8ls_dfxtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.3 0.505 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945 1.125 2.305 1.78 ;
        RECT 1.945 1.78 2.115 2.025 ;
        RECT 1.785 2.025 2.115 2.355 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.705 1.97 9.035 2.98 ;
        RECT 7.805 1.8 9.035 1.97 ;
        RECT 7.805 1.97 8.135 2.98 ;
        RECT 8.865 1.13 9.035 1.8 ;
        RECT 7.82 0.96 9.035 1.13 ;
        RECT 7.82 0.35 8.15 0.96 ;
        RECT 8.7 0.35 9.035 0.96 ;
    END
    ANTENNADIFFAREA 1.116 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
    LAYER li1 ;
      RECT 5.235 1.88 5.405 2.735 ;
      RECT 5.235 1.71 5.86 1.88 ;
      RECT 5.69 1.31 5.86 1.71 ;
      RECT 5.69 1.22 7.13 1.31 ;
      RECT 6.63 1.31 7.13 1.39 ;
      RECT 5.69 1.14 6.8 1.22 ;
      RECT 6.8 1.39 7.13 1.55 ;
      RECT 5.69 0.97 5.86 1.14 ;
      RECT 5.35 0.72 5.86 0.97 ;
      RECT 2.335 2.12 2.505 2.735 ;
      RECT 2.335 1.95 2.645 2.12 ;
      RECT 2.475 1.24 2.645 1.95 ;
      RECT 2.475 1.07 2.995 1.24 ;
      RECT 2.825 0.595 2.995 1.07 ;
      RECT 2.705 2.485 3.035 2.735 ;
      RECT 2.815 2.42 3.035 2.485 ;
      RECT 2.815 2.25 4.385 2.42 ;
      RECT 4.055 1.63 4.385 2.25 ;
      RECT 2.815 1.58 2.985 2.25 ;
      RECT 2.815 1.41 3.345 1.58 ;
      RECT 3.175 0.95 3.345 1.41 ;
      RECT 3.175 0.62 3.535 0.95 ;
      RECT 1.995 2.905 3.375 3.075 ;
      RECT 3.205 2.76 3.375 2.905 ;
      RECT 1.995 2.695 2.165 2.905 ;
      RECT 3.205 2.59 4.385 2.76 ;
      RECT 1.015 2.525 2.165 2.695 ;
      RECT 4.215 2.76 4.385 2.905 ;
      RECT 4.215 2.905 5.955 3.075 ;
      RECT 5.625 2.05 5.955 2.905 ;
      RECT 4.895 1.54 5.065 2.905 ;
      RECT 4.895 1.37 5.52 1.54 ;
      RECT 5.19 1.15 5.52 1.37 ;
      RECT 1.015 2.695 1.475 2.98 ;
      RECT 1.015 1.82 1.475 2.525 ;
      RECT 1.305 1.55 1.475 1.82 ;
      RECT 1.305 1.22 1.765 1.55 ;
      RECT 1.305 0.595 1.475 1.22 ;
      RECT 1.645 0.73 2.655 0.9 ;
      RECT 2.485 0.425 2.655 0.73 ;
      RECT 2.485 0.255 3.875 0.425 ;
      RECT 3.705 0.425 3.875 0.69 ;
      RECT 3.705 0.69 4.68 0.86 ;
      RECT 3.705 0.86 3.875 1.75 ;
      RECT 4.51 0.425 4.68 0.69 ;
      RECT 3.155 1.75 3.875 2.08 ;
      RECT 4.51 0.255 5.995 0.425 ;
      RECT 5.665 0.425 5.995 0.51 ;
      RECT 0.115 2.12 0.445 2.98 ;
      RECT 0.115 1.95 0.845 2.12 ;
      RECT 0.675 1.55 0.845 1.95 ;
      RECT 0.675 1.13 1.135 1.55 ;
      RECT 0.115 0.96 1.135 1.13 ;
      RECT 0.965 0.425 1.135 0.96 ;
      RECT 0.115 0.35 0.445 0.96 ;
      RECT 0.965 0.255 1.815 0.425 ;
      RECT 1.645 0.425 1.815 0.73 ;
      RECT 4.555 1.37 4.725 2.735 ;
      RECT 4.045 1.2 4.725 1.37 ;
      RECT 4.045 1.03 5.02 1.2 ;
      RECT 4.85 0.95 5.02 1.03 ;
      RECT 4.85 0.595 5.18 0.95 ;
      RECT 7.3 1.3 8.665 1.63 ;
      RECT 6.82 1.89 7.15 2.98 ;
      RECT 6.29 1.81 7.47 1.89 ;
      RECT 6.13 1.72 7.47 1.81 ;
      RECT 7.3 1.63 7.47 1.72 ;
      RECT 6.13 1.48 6.46 1.72 ;
      RECT 7.3 1.05 7.47 1.3 ;
      RECT 6.97 0.97 7.47 1.05 ;
      RECT 6.89 0.88 7.47 0.97 ;
      RECT 6.89 0.35 7.14 0.88 ;
      RECT 0 3.245 9.6 3.415 ;
      RECT 9.235 1.82 9.485 3.245 ;
      RECT 3.715 2.93 4.045 3.245 ;
      RECT 6.315 2.45 6.65 3.245 ;
      RECT 7.355 2.06 7.605 3.245 ;
      RECT 0.645 2.29 0.815 3.245 ;
      RECT 1.655 2.865 1.825 3.245 ;
      RECT 8.335 2.14 8.505 3.245 ;
      RECT 0 -0.085 9.6 0.085 ;
      RECT 9.21 0.085 9.46 1.13 ;
      RECT 1.985 0.085 2.315 0.56 ;
      RECT 4.09 0.085 4.34 0.52 ;
      RECT 6.41 0.085 6.66 0.97 ;
      RECT 7.32 0.085 7.65 0.71 ;
      RECT 0.625 0.085 0.795 0.79 ;
      RECT 8.33 0.085 8.5 0.79 ;
  END
END scs8ls_dfxtp_4

MACRO scs8ls_dlclkp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.475 5.155 1.805 ;
    END
    ANTENNAGATEAREA 0.459 ;
  END CLK

  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.47 1.335 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END GATE

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.205 1.55 6.605 2.98 ;
        RECT 6.275 0.35 6.605 1.55 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END GCLK

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.37 2.05 3.775 2.22 ;
      RECT 3.605 1.33 3.775 2.05 ;
      RECT 2.205 1.16 3.775 1.33 ;
      RECT 2.205 1.33 2.535 1.84 ;
      RECT 3.465 0.605 3.775 1.16 ;
      RECT 0.095 0.79 1.215 0.96 ;
      RECT 1.045 0.425 1.215 0.79 ;
      RECT 1.045 0.255 2.955 0.425 ;
      RECT 2.625 0.425 2.955 0.51 ;
      RECT 0.095 1.82 0.445 2.98 ;
      RECT 0.095 1.13 0.265 1.82 ;
      RECT 0.095 0.96 0.445 1.13 ;
      RECT 0.095 0.35 0.445 0.79 ;
      RECT 1.385 2.55 2.285 2.88 ;
      RECT 1.385 2.14 1.555 2.55 ;
      RECT 0.615 1.97 1.555 2.14 ;
      RECT 0.615 1.13 1.555 1.3 ;
      RECT 1.385 0.98 1.555 1.13 ;
      RECT 1.385 0.65 2.26 0.98 ;
      RECT 0.615 1.63 0.785 1.97 ;
      RECT 0.435 1.3 0.785 1.63 ;
      RECT 4.93 2.145 5.26 2.825 ;
      RECT 4.93 1.975 5.535 2.145 ;
      RECT 5.365 1.63 5.535 1.975 ;
      RECT 5.365 1.3 6.035 1.63 ;
      RECT 5.365 1.285 5.615 1.3 ;
      RECT 5.285 0.605 5.615 1.285 ;
      RECT 3.945 2.56 4.26 2.825 ;
      RECT 3.03 2.39 4.26 2.56 ;
      RECT 3.03 2.38 3.2 2.39 ;
      RECT 3.945 1.945 4.26 2.39 ;
      RECT 1.725 2.05 3.2 2.38 ;
      RECT 3.945 1.055 4.205 1.945 ;
      RECT 3.03 1.83 3.2 2.05 ;
      RECT 1.725 1.15 1.995 2.05 ;
      RECT 3.03 1.5 3.435 1.83 ;
      RECT 0 3.245 6.72 3.415 ;
      RECT 2.835 2.73 3.165 3.245 ;
      RECT 0.615 2.31 0.945 3.245 ;
      RECT 4.43 1.975 4.76 3.245 ;
      RECT 5.705 1.945 6.035 3.245 ;
      RECT 0 -0.085 6.72 0.085 ;
      RECT 2.75 0.685 3.295 0.935 ;
      RECT 3.125 0.085 3.295 0.685 ;
      RECT 0.625 0.085 0.875 0.62 ;
      RECT 4.385 0.085 4.715 1.305 ;
      RECT 5.845 0.085 6.095 1.13 ;
    LAYER mcon ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
  END
END scs8ls_dlclkp_1

MACRO scs8ls_dlclkp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.805 0.44 7.135 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END GCLK

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.55 1.445 5.22 1.78 ;
    END
    ANTENNAGATEAREA 0.498 ;
  END CLK

  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.45 1.335 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END GATE

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 4.21 0.575 4.595 1.275 ;
      RECT 4.21 2.075 4.545 2.955 ;
      RECT 4.21 1.885 4.38 2.075 ;
      RECT 3.995 1.555 4.38 1.885 ;
      RECT 4.21 1.275 4.38 1.555 ;
      RECT 5.215 1.95 5.56 2.955 ;
      RECT 5.39 1.61 5.56 1.95 ;
      RECT 5.39 0.94 6.305 1.61 ;
      RECT 5.555 0.575 5.885 0.94 ;
      RECT 3.655 2.1 3.985 2.98 ;
      RECT 3.655 1.385 3.825 2.1 ;
      RECT 2.255 1.215 4.035 1.385 ;
      RECT 2.255 1.385 2.585 1.84 ;
      RECT 3.705 0.605 4.035 1.215 ;
      RECT 0.095 0.77 1.22 0.94 ;
      RECT 1.05 0.425 1.22 0.77 ;
      RECT 1.05 0.255 3.16 0.425 ;
      RECT 2.83 0.425 3.16 0.585 ;
      RECT 0.095 1.82 0.445 2.98 ;
      RECT 0.095 0.94 0.265 1.82 ;
      RECT 0.095 0.35 0.365 0.77 ;
      RECT 2.225 2.22 2.555 2.38 ;
      RECT 1.875 2.05 3.325 2.22 ;
      RECT 3.155 1.885 3.325 2.05 ;
      RECT 1.875 1.45 2.045 2.05 ;
      RECT 3.155 1.555 3.485 1.885 ;
      RECT 1.73 1.12 2.045 1.45 ;
      RECT 1.535 2.55 2.405 2.88 ;
      RECT 1.535 2.12 1.705 2.55 ;
      RECT 0.615 1.95 1.705 2.12 ;
      RECT 0.435 1.11 1.56 1.28 ;
      RECT 1.39 0.95 1.56 1.11 ;
      RECT 1.39 0.62 2.245 0.95 ;
      RECT 0.615 1.55 0.785 1.95 ;
      RECT 0.435 1.28 0.785 1.55 ;
      RECT 0 -0.085 7.68 0.085 ;
      RECT 7.315 0.085 7.565 1.22 ;
      RECT 2.92 0.755 3.535 1.005 ;
      RECT 3.34 0.085 3.535 0.755 ;
      RECT 0.545 0.085 0.88 0.6 ;
      RECT 4.765 0.085 5.095 1.275 ;
      RECT 6.305 0.085 6.635 0.77 ;
      RECT 0 3.245 7.68 3.415 ;
      RECT 7.315 1.82 7.565 3.245 ;
      RECT 2.945 2.65 3.485 3.245 ;
      RECT 0.685 2.29 1.075 3.245 ;
      RECT 4.715 2.075 5.045 3.245 ;
      RECT 5.73 1.95 6.635 3.245 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
  END
END scs8ls_dlclkp_2

MACRO scs8ls_dlclkp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.795 1.55 8.515 1.72 ;
        RECT 7.745 1.72 8.515 1.78 ;
        RECT 6.795 1.72 7.125 2.98 ;
        RECT 7.805 1.38 8.015 1.55 ;
        RECT 7.745 1.78 7.995 2.98 ;
        RECT 6.835 1.21 8.015 1.38 ;
        RECT 6.835 0.35 7.165 1.21 ;
        RECT 7.765 0.35 8.015 1.21 ;
    END
    ANTENNADIFFAREA 1.1032 ;
  END GCLK

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.4 1.36 5.07 1.78 ;
    END
    ANTENNAGATEAREA 0.516 ;
  END CLK

  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.53 1.43 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END GATE

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 4.28 0.515 4.61 0.85 ;
      RECT 3.815 0.255 4.61 0.515 ;
      RECT 3.645 2.18 3.995 2.35 ;
      RECT 3.825 1.61 3.995 2.18 ;
      RECT 3.825 1.53 4.155 1.61 ;
      RECT 2.305 1.36 4.155 1.53 ;
      RECT 2.305 1.53 2.635 1.805 ;
      RECT 5.24 1.99 5.57 2.98 ;
      RECT 5.24 1.82 6.35 1.99 ;
      RECT 5.975 1.13 6.35 1.82 ;
      RECT 5.6 0.67 6.35 1.13 ;
      RECT 5.6 0.35 5.975 0.67 ;
      RECT 2.815 1.02 5.43 1.19 ;
      RECT 5.26 1.19 5.43 1.3 ;
      RECT 5.26 1.3 5.805 1.63 ;
      RECT 0.115 0.85 1.265 1.02 ;
      RECT 1.095 0.425 1.265 0.85 ;
      RECT 1.095 0.255 3.145 0.425 ;
      RECT 2.815 0.425 3.145 1.02 ;
      RECT 0.115 1.82 0.54 2.98 ;
      RECT 0.115 1.02 0.365 1.82 ;
      RECT 0.115 0.35 0.365 0.85 ;
      RECT 4.205 2.69 4.535 2.97 ;
      RECT 3.305 2.52 4.535 2.69 ;
      RECT 4.205 2.09 4.535 2.52 ;
      RECT 3.305 2.35 3.475 2.52 ;
      RECT 1.775 2.05 3.475 2.35 ;
      RECT 3.305 1.96 3.475 2.05 ;
      RECT 1.775 1.15 2.065 2.05 ;
      RECT 3.305 1.7 3.655 1.96 ;
      RECT 1.435 2.52 2.485 2.85 ;
      RECT 1.435 2.14 1.605 2.52 ;
      RECT 0.71 1.97 1.605 2.14 ;
      RECT 0.535 1.19 1.605 1.36 ;
      RECT 1.435 0.98 1.605 1.19 ;
      RECT 1.435 0.65 2.33 0.98 ;
      RECT 0.71 1.55 0.88 1.97 ;
      RECT 0.535 1.36 0.88 1.55 ;
      RECT 0 -0.085 8.64 0.085 ;
      RECT 8.195 0.085 8.525 1.04 ;
      RECT 0.55 0.085 0.925 0.68 ;
      RECT 3.315 0.085 3.645 0.85 ;
      RECT 4.78 0.085 5.11 0.85 ;
      RECT 6.16 0.085 6.655 0.5 ;
      RECT 7.335 0.085 7.585 1.04 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 8.195 1.95 8.525 3.245 ;
      RECT 3.11 2.86 3.44 3.245 ;
      RECT 0.785 2.31 1.16 3.245 ;
      RECT 5.74 2.16 6.625 3.245 ;
      RECT 4.74 2.09 5.07 3.245 ;
      RECT 7.295 1.89 7.545 3.245 ;
    LAYER mcon ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
  END
END scs8ls_dlclkp_4

MACRO scs8ls_dlrbn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.26 0.835 1.9 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END D

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.875 1.18 6.18 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END RESETB

  PIN GATEN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.26 1.335 1.9 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END GATEN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.565 0.35 7.115 1.05 ;
        RECT 6.945 1.05 7.115 1.72 ;
        RECT 6.69 1.72 7.115 2.85 ;
    END
    ANTENNADIFFAREA 0.5357 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.195 1.82 8.53 2.98 ;
        RECT 8.36 1.13 8.53 1.82 ;
        RECT 8.245 0.35 8.53 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END QN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.12 2.905 4.29 3.075 ;
      RECT 3.12 2.14 3.29 2.905 ;
      RECT 3.96 2.05 4.29 2.905 ;
      RECT 3.12 1.97 3.45 2.14 ;
      RECT 3.28 1.45 3.45 1.97 ;
      RECT 3.28 1.3 3.61 1.45 ;
      RECT 2.185 1.13 3.61 1.3 ;
      RECT 2.185 1.3 2.555 1.55 ;
      RECT 3.28 1.12 3.61 1.13 ;
      RECT 2.385 1.55 2.555 2.22 ;
      RECT 1.405 2.22 2.555 2.39 ;
      RECT 1.405 2.39 1.675 2.56 ;
      RECT 1.405 2.1 1.675 2.22 ;
      RECT 1.505 1.09 1.675 2.1 ;
      RECT 1.13 0.35 1.675 1.09 ;
      RECT 1.845 1.72 2.215 2.05 ;
      RECT 1.845 0.96 2.015 1.72 ;
      RECT 1.845 0.95 2.175 0.96 ;
      RECT 1.845 0.78 4.205 0.95 ;
      RECT 3.875 0.95 4.205 1.45 ;
      RECT 1.845 0.35 2.175 0.78 ;
      RECT 3.46 2.405 3.79 2.735 ;
      RECT 3.62 1.79 3.79 2.405 ;
      RECT 3.62 1.62 4.725 1.79 ;
      RECT 4.375 1.55 4.725 1.62 ;
      RECT 4.375 1.22 5.12 1.55 ;
      RECT 4.375 0.61 4.545 1.22 ;
      RECT 3.405 0.36 4.545 0.61 ;
      RECT 1.065 2.73 2.015 2.9 ;
      RECT 1.845 2.56 2.91 2.73 ;
      RECT 1.065 2.24 1.235 2.73 ;
      RECT 2.74 1.8 2.91 2.56 ;
      RECT 0.095 2.07 1.235 2.24 ;
      RECT 2.74 1.47 3.07 1.8 ;
      RECT 0.095 0.54 0.45 1.09 ;
      RECT 0.095 2.24 0.365 2.98 ;
      RECT 0.095 1.09 0.265 2.07 ;
      RECT 6.35 1.22 6.775 1.55 ;
      RECT 5.615 2.29 5.945 2.85 ;
      RECT 4.53 1.96 5.945 2.29 ;
      RECT 5.29 1.89 5.945 1.96 ;
      RECT 5.29 1.72 6.52 1.89 ;
      RECT 6.35 1.55 6.52 1.72 ;
      RECT 5.29 1.05 5.46 1.72 ;
      RECT 5.21 0.35 5.46 1.05 ;
      RECT 7.285 1.63 7.535 2.78 ;
      RECT 7.285 1.3 8.19 1.63 ;
      RECT 7.285 0.54 7.56 1.3 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 7.745 1.82 8.01 3.245 ;
      RECT 2.505 2.9 2.835 3.245 ;
      RECT 4.68 2.52 5.445 3.245 ;
      RECT 6.115 2.06 6.445 3.245 ;
      RECT 0.565 2.41 0.895 3.245 ;
      RECT 0 -0.085 8.64 0.085 ;
      RECT 7.745 0.085 8.075 1.13 ;
      RECT 0.63 0.085 0.96 1.09 ;
      RECT 2.345 0.085 2.915 0.6 ;
      RECT 4.73 0.085 4.98 1.03 ;
      RECT 6.03 0.085 6.36 1.01 ;
    LAYER mcon ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
  END
END scs8ls_dlrbn_1

MACRO scs8ls_dlrbn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.225 1.82 8.575 2.98 ;
        RECT 8.405 1.05 8.575 1.82 ;
        RECT 8.205 0.88 8.575 1.05 ;
    END
    ANTENNADIFFAREA 0.5728 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.285 0.77 6.615 1.13 ;
        RECT 6.285 1.13 6.455 1.82 ;
        RECT 6.26 1.82 6.59 2.07 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END Q

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.57 1.18 6.115 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END RESETB

  PIN GATEN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.975 1.26 1.285 1.93 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END GATEN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.26 0.805 1.93 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.985 2.65 1.965 2.82 ;
      RECT 1.795 2.48 2.83 2.65 ;
      RECT 0.985 2.27 1.155 2.65 ;
      RECT 2.66 1.8 2.83 2.48 ;
      RECT 0.085 2.1 1.155 2.27 ;
      RECT 2.66 1.47 2.985 1.8 ;
      RECT 0.085 2.27 0.445 2.98 ;
      RECT 0.085 0.54 0.445 1.09 ;
      RECT 0.085 1.09 0.255 2.1 ;
      RECT 3.01 2.905 4.165 3.075 ;
      RECT 3.01 2.14 3.18 2.905 ;
      RECT 3.835 2.05 4.165 2.905 ;
      RECT 3.01 1.97 3.325 2.14 ;
      RECT 3.155 1.45 3.325 1.97 ;
      RECT 3.155 1.3 3.53 1.45 ;
      RECT 2.135 1.13 3.53 1.3 ;
      RECT 2.135 1.3 2.475 1.55 ;
      RECT 3.155 1.12 3.53 1.13 ;
      RECT 2.305 1.55 2.475 2.14 ;
      RECT 1.325 2.14 2.475 2.31 ;
      RECT 1.325 2.31 1.625 2.48 ;
      RECT 1.325 2.1 1.625 2.14 ;
      RECT 1.455 1.09 1.625 2.1 ;
      RECT 1.125 0.35 1.625 1.09 ;
      RECT 1.795 1.72 2.135 1.97 ;
      RECT 1.795 0.96 1.965 1.72 ;
      RECT 1.795 0.95 2.125 0.96 ;
      RECT 1.795 0.78 3.885 0.95 ;
      RECT 3.715 0.95 3.885 1.225 ;
      RECT 1.795 0.35 2.125 0.78 ;
      RECT 3.715 1.225 4.13 1.54 ;
      RECT 7.215 1.22 8.23 1.55 ;
      RECT 7.215 1.55 7.545 2.86 ;
      RECT 7.215 0.35 7.545 1.22 ;
      RECT 5.31 2.35 6.955 2.41 ;
      RECT 4.375 2.24 6.955 2.35 ;
      RECT 6.785 1.65 6.955 2.24 ;
      RECT 6.625 1.32 6.955 1.65 ;
      RECT 5.31 2.41 5.64 2.98 ;
      RECT 4.375 2.05 5.64 2.24 ;
      RECT 5.23 1.82 5.64 2.05 ;
      RECT 5.23 1.13 5.4 1.82 ;
      RECT 4.875 0.35 5.4 1.13 ;
      RECT 3.35 2.405 3.665 2.735 ;
      RECT 3.495 1.88 3.665 2.405 ;
      RECT 3.495 1.71 5.06 1.88 ;
      RECT 4.735 1.35 5.06 1.71 ;
      RECT 4.3 1.055 4.47 1.71 ;
      RECT 4.055 0.885 4.47 1.055 ;
      RECT 4.055 0.61 4.225 0.885 ;
      RECT 3.325 0.36 4.225 0.61 ;
      RECT 0 -0.085 9.12 0.085 ;
      RECT 8.745 0.085 9.005 1.13 ;
      RECT 6.785 0.085 7.045 1.05 ;
      RECT 7.775 0.085 8.035 1.05 ;
      RECT 0.625 0.085 0.955 1.09 ;
      RECT 2.295 0.085 2.835 0.6 ;
      RECT 4.395 0.085 4.645 0.715 ;
      RECT 5.695 0.085 6.025 1.01 ;
      RECT 0 3.245 9.12 3.415 ;
      RECT 8.755 1.82 9.005 3.245 ;
      RECT 6.71 2.58 7.04 3.245 ;
      RECT 7.775 1.82 8.025 3.245 ;
      RECT 2.425 2.82 2.755 3.245 ;
      RECT 4.525 2.65 5.14 3.245 ;
      RECT 5.81 2.58 6.14 3.245 ;
      RECT 0.645 2.44 0.815 3.245 ;
    LAYER mcon ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
  END
END scs8ls_dlrbn_2

MACRO scs8ls_dlrbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.425 1.18 5.795 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END RESETB

  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.975 1.45 1.305 1.78 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END GATE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.2 2.06 6.67 2.98 ;
        RECT 6.5 1.18 6.67 2.06 ;
        RECT 6.13 1.01 6.67 1.18 ;
        RECT 6.13 0.35 6.46 1.01 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.71 0.35 8.055 1.04 ;
        RECT 7.885 1.04 8.055 1.82 ;
        RECT 7.715 1.82 8.055 2.98 ;
    END
    ANTENNADIFFAREA 0.6042 ;
  END QN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.45 0.805 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.185 1.97 1.645 2.22 ;
      RECT 1.475 1.75 1.645 1.97 ;
      RECT 1.475 1.42 1.875 1.75 ;
      RECT 1.475 1.28 1.645 1.42 ;
      RECT 1.185 0.75 1.645 1.28 ;
      RECT 1.185 0.58 2.99 0.75 ;
      RECT 2.82 0.51 2.99 0.58 ;
      RECT 1.185 0.5 1.645 0.58 ;
      RECT 2.82 0.255 3.905 0.51 ;
      RECT 2.855 2.905 4.015 3.075 ;
      RECT 2.855 2.14 3.025 2.905 ;
      RECT 3.685 2.05 4.015 2.905 ;
      RECT 2.855 1.97 3.175 2.14 ;
      RECT 3.005 1.48 3.175 1.97 ;
      RECT 3.005 1.3 3.395 1.48 ;
      RECT 2.045 1.25 3.395 1.3 ;
      RECT 2.045 1.3 2.215 1.94 ;
      RECT 1.825 1.13 3.395 1.25 ;
      RECT 1.815 1.94 2.215 2.22 ;
      RECT 1.825 0.92 2.215 1.13 ;
      RECT 3.195 2.405 3.515 2.735 ;
      RECT 3.345 1.82 3.515 2.405 ;
      RECT 3.345 1.65 4.915 1.82 ;
      RECT 4.585 1.35 4.915 1.65 ;
      RECT 3.58 0.96 3.75 1.65 ;
      RECT 3.19 0.71 3.75 0.96 ;
      RECT 0.095 2.39 2.675 2.56 ;
      RECT 2.505 1.8 2.675 2.39 ;
      RECT 2.505 1.47 2.835 1.8 ;
      RECT 0.095 2.56 0.445 2.85 ;
      RECT 0.095 1.97 0.445 2.39 ;
      RECT 0.095 0.69 0.445 1.28 ;
      RECT 0.095 1.28 0.265 1.97 ;
      RECT 6.84 1.32 7.715 1.65 ;
      RECT 6.84 1.65 7.01 2.98 ;
      RECT 6.84 0.84 7.02 1.32 ;
      RECT 6.69 0.35 7.02 0.84 ;
      RECT 5.085 1.72 6.33 1.89 ;
      RECT 6.005 1.35 6.33 1.72 ;
      RECT 5.25 2.32 5.58 2.98 ;
      RECT 4.225 1.99 5.58 2.32 ;
      RECT 5.085 1.89 5.58 1.99 ;
      RECT 5.085 1.13 5.255 1.72 ;
      RECT 4.8 0.35 5.255 1.13 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 7.21 2.1 7.54 3.245 ;
      RECT 0.65 2.73 0.98 3.245 ;
      RECT 2.35 2.73 2.685 3.245 ;
      RECT 4.405 2.65 5.08 3.245 ;
      RECT 5.78 2.06 6.03 3.245 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 7.2 0.085 7.53 0.94 ;
      RECT 5.62 0.085 5.95 1.01 ;
      RECT 0.625 0.085 0.955 1.28 ;
      RECT 2.32 0.085 2.65 0.41 ;
      RECT 4.24 0.085 4.57 1.06 ;
    LAYER mcon ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
  END
END scs8ls_dlrbp_1

MACRO scs8ls_dlrbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845 1.13 7.075 1.8 ;
        RECT 6.295 1.8 7.075 1.97 ;
        RECT 6.15 0.96 7.075 1.13 ;
        RECT 6.295 1.97 6.465 2.98 ;
        RECT 6.15 0.35 6.48 0.96 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.225 1.82 8.585 2.98 ;
        RECT 8.415 1.13 8.585 1.82 ;
        RECT 8.245 0.35 8.585 1.13 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END QN

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.435 1.18 5.785 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END RESETB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.45 0.805 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END D

  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.975 1.18 1.285 1.55 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END GATE

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.315 1.82 3.485 2.735 ;
      RECT 3.315 1.65 4.925 1.82 ;
      RECT 4.605 1.35 4.925 1.65 ;
      RECT 3.57 0.96 3.74 1.65 ;
      RECT 3.18 0.79 3.74 0.96 ;
      RECT 0.085 2.36 2.805 2.53 ;
      RECT 2.485 1.47 2.805 2.36 ;
      RECT 0.085 2.53 0.445 2.82 ;
      RECT 0.085 1.95 0.445 2.36 ;
      RECT 0.085 0.54 0.445 1.13 ;
      RECT 0.085 1.13 0.255 1.95 ;
      RECT 5.955 1.3 6.65 1.63 ;
      RECT 5.235 2.32 5.565 2.98 ;
      RECT 4.245 1.99 5.565 2.32 ;
      RECT 5.095 1.89 5.565 1.99 ;
      RECT 5.095 1.72 6.125 1.89 ;
      RECT 5.955 1.63 6.125 1.72 ;
      RECT 5.095 1.13 5.265 1.72 ;
      RECT 4.79 0.35 5.265 1.13 ;
      RECT 2.975 2.905 4.035 3.075 ;
      RECT 3.705 2.05 4.035 2.905 ;
      RECT 2.975 1.48 3.145 2.905 ;
      RECT 2.975 1.3 3.385 1.48 ;
      RECT 2.035 1.17 3.385 1.3 ;
      RECT 2.035 1.3 2.205 1.94 ;
      RECT 1.795 1.13 3.385 1.17 ;
      RECT 1.795 1.94 2.205 2.19 ;
      RECT 1.795 0.92 2.205 1.13 ;
      RECT 1.185 1.94 1.625 2.19 ;
      RECT 1.455 1.67 1.625 1.94 ;
      RECT 1.455 1.34 1.865 1.67 ;
      RECT 1.455 1.01 1.625 1.34 ;
      RECT 1.125 0.75 1.625 1.01 ;
      RECT 1.125 0.58 2.98 0.75 ;
      RECT 2.81 0.51 2.98 0.58 ;
      RECT 1.125 0.35 1.625 0.58 ;
      RECT 2.81 0.255 3.895 0.51 ;
      RECT 7.245 1.3 8.245 1.63 ;
      RECT 7.245 1.63 7.555 2.86 ;
      RECT 7.245 1.13 7.555 1.3 ;
      RECT 7.245 0.45 7.575 1.13 ;
      RECT 0 -0.085 9.12 0.085 ;
      RECT 8.755 0.085 9.005 1.13 ;
      RECT 6.65 0.085 6.98 0.79 ;
      RECT 7.745 0.085 8.075 1.13 ;
      RECT 0.625 0.085 0.955 1.01 ;
      RECT 2.305 0.085 2.64 0.41 ;
      RECT 4.23 0.085 4.56 1.06 ;
      RECT 5.61 0.085 5.94 1.01 ;
      RECT 0 3.245 9.12 3.415 ;
      RECT 8.755 1.82 9.005 3.245 ;
      RECT 6.665 2.14 6.995 3.245 ;
      RECT 7.725 1.82 8.055 3.245 ;
      RECT 0.65 2.7 0.98 3.245 ;
      RECT 2.33 2.7 2.695 3.245 ;
      RECT 4.425 2.65 5.065 3.245 ;
      RECT 5.735 2.06 6.065 3.245 ;
    LAYER mcon ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_dlrbp_2

MACRO scs8ls_dlrtn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.755 1.82 7.115 2.98 ;
        RECT 6.945 1.13 7.115 1.82 ;
        RECT 6.73 0.35 7.115 1.13 ;
    END
    ANTENNADIFFAREA 0.6005 ;
  END Q

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.18 6.235 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END RESETB

  PIN GATEN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.45 1.335 1.78 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END GATEN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.45 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 6.415 1.32 6.775 1.65 ;
      RECT 5.635 2.36 5.965 2.86 ;
      RECT 4.485 2.03 5.965 2.36 ;
      RECT 5.465 1.89 5.965 2.03 ;
      RECT 5.465 1.72 6.585 1.89 ;
      RECT 6.415 1.65 6.585 1.72 ;
      RECT 5.465 1.13 5.635 1.72 ;
      RECT 5.24 0.35 5.635 1.13 ;
      RECT 0.095 0.58 2.865 0.75 ;
      RECT 2.535 0.75 2.865 1.59 ;
      RECT 0.095 1.95 0.45 2.83 ;
      RECT 0.095 0.75 0.445 1.25 ;
      RECT 0.095 1.25 0.265 1.95 ;
      RECT 3.255 2.18 3.745 2.35 ;
      RECT 3.575 1.86 3.745 2.18 ;
      RECT 3.575 1.69 5.07 1.86 ;
      RECT 4.9 1.63 5.07 1.69 ;
      RECT 4.9 1.3 5.295 1.63 ;
      RECT 4.9 1.02 5.07 1.3 ;
      RECT 3.815 0.85 5.07 1.02 ;
      RECT 3.815 0.35 4.145 0.85 ;
      RECT 1.845 2.01 2.245 2.35 ;
      RECT 1.845 1.84 3.405 2.01 ;
      RECT 3.075 1.52 3.405 1.84 ;
      RECT 2.075 1.17 2.245 1.84 ;
      RECT 3.075 1.19 4.335 1.52 ;
      RECT 1.845 0.92 2.245 1.17 ;
      RECT 1.19 2.69 1.675 2.83 ;
      RECT 1.19 2.52 4.245 2.69 ;
      RECT 3.915 2.03 4.245 2.52 ;
      RECT 1.19 1.95 1.675 2.52 ;
      RECT 1.505 1.67 1.675 1.95 ;
      RECT 1.505 1.34 1.905 1.67 ;
      RECT 1.505 1.25 1.675 1.34 ;
      RECT 1.065 0.92 1.675 1.25 ;
      RECT 0 -0.085 7.2 0.085 ;
      RECT 0.625 0.085 0.955 0.41 ;
      RECT 2.355 0.085 3.2 0.41 ;
      RECT 4.67 0.085 5.01 0.68 ;
      RECT 6.14 0.085 6.47 1.01 ;
      RECT 0 3.245 7.2 3.415 ;
      RECT 2.3 2.86 2.63 3.245 ;
      RECT 4.635 2.53 5.43 3.245 ;
      RECT 6.255 2.06 6.585 3.245 ;
      RECT 0.655 1.95 0.985 3.245 ;
    LAYER mcon ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
  END
END scs8ls_dlrtn_1

MACRO scs8ls_dlrtn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845 1.82 7.535 2.98 ;
        RECT 7.365 1.47 7.535 1.82 ;
        RECT 7.205 0.35 7.535 1.47 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END Q

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.18 6.305 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END RESETB

  PIN GATEN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.45 1.335 1.78 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END GATEN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.45 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.335 2.18 3.825 2.35 ;
      RECT 3.655 1.86 3.825 2.18 ;
      RECT 3.655 1.69 5.375 1.86 ;
      RECT 4.97 1.35 5.375 1.69 ;
      RECT 4.97 1.02 5.14 1.35 ;
      RECT 3.895 0.85 5.14 1.02 ;
      RECT 3.895 0.35 4.225 0.85 ;
      RECT 1.845 2.01 2.245 2.35 ;
      RECT 1.845 1.84 3.485 2.01 ;
      RECT 3.155 1.52 3.485 1.84 ;
      RECT 2.075 1.17 2.245 1.84 ;
      RECT 3.155 1.19 4.415 1.52 ;
      RECT 1.845 0.92 2.245 1.17 ;
      RECT 0.095 0.58 2.945 0.75 ;
      RECT 2.615 0.75 2.945 1.59 ;
      RECT 0.095 1.95 0.615 2.83 ;
      RECT 0.095 0.75 0.445 1.25 ;
      RECT 0.095 1.25 0.265 1.95 ;
      RECT 1.285 2.69 1.675 2.83 ;
      RECT 1.285 2.52 4.325 2.69 ;
      RECT 3.995 2.03 4.325 2.52 ;
      RECT 1.285 1.95 1.675 2.52 ;
      RECT 1.505 1.67 1.675 1.95 ;
      RECT 1.505 1.34 1.905 1.67 ;
      RECT 1.505 1.25 1.675 1.34 ;
      RECT 1.135 0.92 1.675 1.25 ;
      RECT 5.715 2.36 6.045 2.98 ;
      RECT 4.565 2.03 6.045 2.36 ;
      RECT 5.545 1.89 6.045 2.03 ;
      RECT 5.545 1.72 6.675 1.89 ;
      RECT 6.505 1.65 6.675 1.72 ;
      RECT 6.505 1.32 6.845 1.65 ;
      RECT 5.545 1.13 5.715 1.72 ;
      RECT 5.31 0.35 5.715 1.13 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 7.705 0.085 8.035 1.13 ;
      RECT 0.625 0.085 0.955 0.41 ;
      RECT 2.38 0.085 3.28 0.41 ;
      RECT 4.75 0.085 5.08 0.68 ;
      RECT 6.13 0.085 7.035 1.01 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 7.705 1.82 8.045 3.245 ;
      RECT 2.38 2.86 2.71 3.245 ;
      RECT 4.715 2.63 5.545 3.245 ;
      RECT 6.32 2.06 6.65 3.245 ;
      RECT 0.785 1.95 1.115 3.245 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
  END
END scs8ls_dlrtn_2

MACRO scs8ls_dlrtn_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.795 0.8 9.475 0.96 ;
        RECT 7.935 0.96 9.475 1.13 ;
        RECT 8.795 0.36 8.985 0.8 ;
        RECT 9.245 1.13 9.475 1.8 ;
        RECT 7.935 0.36 8.125 0.96 ;
        RECT 8.545 1.8 9.475 1.96 ;
        RECT 7.545 1.96 9.475 1.97 ;
        RECT 7.545 1.97 8.875 2.13 ;
        RECT 7.545 2.13 7.875 2.98 ;
        RECT 8.545 2.13 8.875 2.98 ;
    END
    ANTENNADIFFAREA 1.1984 ;
  END Q

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.32 1.12 7.555 1.45 ;
    END
    ANTENNAGATEAREA 0.444 ;
  END RESETB

  PIN GATEN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.975 1.45 1.29 1.78 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END GATEN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.45 0.805 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 5.155 0.425 5.485 0.95 ;
      RECT 5.155 0.255 6.265 0.425 ;
      RECT 6.015 0.425 6.265 0.77 ;
      RECT 6.015 0.77 7.205 0.95 ;
      RECT 6.945 0.355 7.205 0.77 ;
      RECT 1.8 2.09 2.205 2.43 ;
      RECT 1.8 1.92 3.36 2.09 ;
      RECT 3.03 1.52 3.36 1.92 ;
      RECT 2.035 1.25 2.205 1.92 ;
      RECT 3.03 1.19 4.26 1.52 ;
      RECT 1.8 1 2.205 1.25 ;
      RECT 0.085 0.66 2.82 0.83 ;
      RECT 2.49 0.83 2.82 1.67 ;
      RECT 0.085 1.95 0.475 2.83 ;
      RECT 0.085 0.83 0.445 1.25 ;
      RECT 0.085 1.25 0.255 1.95 ;
      RECT 1.145 2.77 1.63 2.83 ;
      RECT 1.145 2.6 4.2 2.77 ;
      RECT 3.87 2.03 4.2 2.6 ;
      RECT 1.145 1.95 1.63 2.6 ;
      RECT 1.46 1.75 1.63 1.95 ;
      RECT 1.46 1.42 1.865 1.75 ;
      RECT 1.46 1.25 1.63 1.42 ;
      RECT 1.135 1 1.63 1.25 ;
      RECT 3.18 2.26 3.7 2.43 ;
      RECT 3.53 1.86 3.7 2.26 ;
      RECT 3.53 1.69 5.22 1.86 ;
      RECT 4.815 1.12 5.22 1.69 ;
      RECT 4.815 1.02 4.985 1.12 ;
      RECT 3.74 0.85 4.985 1.02 ;
      RECT 3.74 0.4 4.07 0.85 ;
      RECT 5.49 1.62 9.075 1.63 ;
      RECT 7.725 1.3 9.075 1.62 ;
      RECT 6.49 1.79 6.82 2.96 ;
      RECT 5.49 1.63 7.895 1.79 ;
      RECT 5.49 2.36 5.82 2.96 ;
      RECT 4.44 2.03 5.82 2.36 ;
      RECT 5.49 1.79 5.82 2.03 ;
      RECT 5.665 0.595 5.835 1.62 ;
      RECT 0 -0.085 9.6 0.085 ;
      RECT 9.155 0.085 9.485 0.63 ;
      RECT 0.625 0.085 0.955 0.49 ;
      RECT 2.31 0.085 3.125 0.49 ;
      RECT 4.595 0.085 4.925 0.68 ;
      RECT 6.445 0.085 6.775 0.6 ;
      RECT 7.435 0.085 7.765 0.95 ;
      RECT 8.295 0.085 8.625 0.79 ;
      RECT 0 3.245 9.6 3.415 ;
      RECT 9.045 2.14 9.375 3.245 ;
      RECT 2.255 2.94 2.585 3.245 ;
      RECT 4.59 2.63 5.32 3.245 ;
      RECT 5.99 2.08 6.32 3.245 ;
      RECT 7.045 2.08 7.375 3.245 ;
      RECT 0.645 1.95 0.975 3.245 ;
      RECT 8.045 2.3 8.375 3.245 ;
    LAYER mcon ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
  END
END scs8ls_dlrtn_4

MACRO scs8ls_dlrtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.3 0.375 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END D

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.435 1.35 5.765 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END RESETB

  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.93 1.45 1.285 1.78 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END GATE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.1 0.35 6.635 0.84 ;
        RECT 6.465 0.84 6.635 1.82 ;
        RECT 6.275 1.82 6.635 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.905 2.905 4.045 3.075 ;
      RECT 2.905 2.14 3.075 2.905 ;
      RECT 3.715 2.065 4.045 2.905 ;
      RECT 2.905 1.97 3.195 2.14 ;
      RECT 3.025 1.45 3.195 1.97 ;
      RECT 3.025 1.28 3.325 1.45 ;
      RECT 1.795 1.11 3.325 1.28 ;
      RECT 2 1.28 2.17 2.02 ;
      RECT 1.795 2.02 2.17 2.22 ;
      RECT 3.245 2.405 3.535 2.735 ;
      RECT 3.365 1.895 3.535 2.405 ;
      RECT 3.365 1.725 4.925 1.895 ;
      RECT 4.665 1.47 4.925 1.725 ;
      RECT 3.495 0.925 3.665 1.725 ;
      RECT 3.19 0.595 3.665 0.925 ;
      RECT 1.15 1.97 1.625 2.22 ;
      RECT 1.455 1.78 1.625 1.97 ;
      RECT 1.455 1.45 1.83 1.78 ;
      RECT 1.455 1.13 1.625 1.45 ;
      RECT 1.235 0.94 1.625 1.13 ;
      RECT 1.235 0.77 3.02 0.94 ;
      RECT 2.85 0.425 3.02 0.77 ;
      RECT 1.235 0.35 1.625 0.77 ;
      RECT 2.85 0.255 4.005 0.425 ;
      RECT 3.835 0.425 4.005 1.225 ;
      RECT 3.835 1.225 4.095 1.555 ;
      RECT 0.115 2.39 2.695 2.56 ;
      RECT 2.525 1.8 2.695 2.39 ;
      RECT 2.525 1.47 2.855 1.8 ;
      RECT 0.115 2.56 0.445 2.98 ;
      RECT 0.115 2.1 0.715 2.39 ;
      RECT 0.545 1.13 0.715 2.1 ;
      RECT 0.22 0.54 0.715 1.13 ;
      RECT 4.77 1.01 6.295 1.18 ;
      RECT 5.975 1.18 6.295 1.55 ;
      RECT 5.245 2.38 5.575 2.98 ;
      RECT 4.305 2.065 5.575 2.38 ;
      RECT 5.095 1.95 5.575 2.065 ;
      RECT 5.095 1.18 5.265 1.95 ;
      RECT 4.77 0.35 5.1 1.01 ;
      RECT 0 3.245 6.72 3.415 ;
      RECT 0.615 2.73 0.945 3.245 ;
      RECT 2.33 2.73 2.705 3.245 ;
      RECT 4.435 2.65 5.075 3.245 ;
      RECT 5.745 1.95 6.075 3.245 ;
      RECT 0 -0.085 6.72 0.085 ;
      RECT 0.885 0.085 1.055 1.13 ;
      RECT 2.295 0.085 2.68 0.6 ;
      RECT 4.21 0.085 4.54 0.81 ;
      RECT 5.59 0.085 5.92 0.84 ;
    LAYER mcon ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
  END
END scs8ls_dlrtp_1

MACRO scs8ls_dlrtp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845 1.13 7.075 1.8 ;
        RECT 6.415 1.8 7.075 1.97 ;
        RECT 6.255 0.96 7.075 1.13 ;
        RECT 6.415 1.97 6.585 2.06 ;
        RECT 6.255 0.35 6.585 0.96 ;
        RECT 6.255 2.06 6.585 2.98 ;
    END
    ANTENNADIFFAREA 0.5674 ;
  END Q

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.435 1.18 5.84 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END RESETB

  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.18 1.285 1.55 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END GATE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.45 0.515 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 6.05 1.3 6.675 1.63 ;
      RECT 5.255 2.38 5.585 2.98 ;
      RECT 4.3 2.1 5.585 2.38 ;
      RECT 5.095 1.89 5.585 2.1 ;
      RECT 5.095 1.72 6.22 1.89 ;
      RECT 6.05 1.63 6.22 1.72 ;
      RECT 5.095 1.13 5.265 1.72 ;
      RECT 4.845 0.35 5.265 1.13 ;
      RECT 0.115 2.44 2.68 2.61 ;
      RECT 2.51 1.77 2.68 2.44 ;
      RECT 2.51 1.44 2.84 1.77 ;
      RECT 0.115 2.61 0.445 2.82 ;
      RECT 0.115 1.95 0.855 2.44 ;
      RECT 0.685 1.28 0.855 1.95 ;
      RECT 0.14 1.11 0.855 1.28 ;
      RECT 0.14 0.54 0.47 1.11 ;
      RECT 3.23 2.405 3.56 2.735 ;
      RECT 3.39 1.93 3.56 2.405 ;
      RECT 3.39 1.76 4.925 1.93 ;
      RECT 4.66 1.35 4.925 1.76 ;
      RECT 3.485 0.845 3.655 1.76 ;
      RECT 3.205 0.595 3.715 0.845 ;
      RECT 2.89 2.905 4.06 3.075 ;
      RECT 2.89 2.11 3.06 2.905 ;
      RECT 3.73 2.1 4.06 2.905 ;
      RECT 2.89 1.94 3.22 2.11 ;
      RECT 3.05 1.45 3.22 1.94 ;
      RECT 3.05 1.25 3.315 1.45 ;
      RECT 1.795 1.08 3.315 1.25 ;
      RECT 2.06 1.25 2.23 1.94 ;
      RECT 1.795 0.92 2.23 1.08 ;
      RECT 1.825 1.94 2.23 2.27 ;
      RECT 1.185 1.94 1.625 2.27 ;
      RECT 1.455 1.75 1.625 1.94 ;
      RECT 1.455 1.42 1.89 1.75 ;
      RECT 1.455 1.01 1.625 1.42 ;
      RECT 1.15 0.75 1.625 1.01 ;
      RECT 1.15 0.58 2.975 0.75 ;
      RECT 2.805 0.425 2.975 0.58 ;
      RECT 1.15 0.35 1.625 0.58 ;
      RECT 2.805 0.255 4.09 0.425 ;
      RECT 3.92 0.425 4.09 1.26 ;
      RECT 3.825 1.26 4.09 1.59 ;
      RECT 0 -0.085 7.2 0.085 ;
      RECT 6.755 0.085 7.085 0.79 ;
      RECT 0.65 0.085 0.98 0.94 ;
      RECT 2.305 0.085 2.635 0.41 ;
      RECT 4.285 0.085 4.615 0.845 ;
      RECT 5.755 0.085 6.085 1.01 ;
      RECT 0 3.245 7.2 3.415 ;
      RECT 6.755 2.14 7.085 3.245 ;
      RECT 0.65 2.78 0.98 3.245 ;
      RECT 2.28 2.78 2.61 3.245 ;
      RECT 4.45 2.65 5.085 3.245 ;
      RECT 5.755 2.06 6.085 3.245 ;
    LAYER mcon ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
  END
END scs8ls_dlrtp_2

MACRO scs8ls_dlrtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.765 1.13 8.995 1.8 ;
        RECT 7.175 1.8 8.995 1.97 ;
        RECT 7.385 0.88 8.995 1.13 ;
        RECT 7.175 1.97 7.425 2.98 ;
        RECT 8.095 1.97 8.425 2.98 ;
        RECT 7.385 0.365 7.645 0.88 ;
        RECT 8.315 0.365 8.505 0.88 ;
    END
    ANTENNADIFFAREA 1.1648 ;
  END Q

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.12 6.595 1.45 ;
    END
    ANTENNAGATEAREA 0.444 ;
  END RESETB

  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.45 1.29 1.78 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END GATE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.45 0.515 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 4.67 0.45 5 1.03 ;
      RECT 4.67 0.28 5.785 0.45 ;
      RECT 5.535 0.45 5.785 0.77 ;
      RECT 5.535 0.77 6.725 0.95 ;
      RECT 6.465 0.345 6.725 0.77 ;
      RECT 3.185 2.405 3.465 2.735 ;
      RECT 3.295 1.895 3.465 2.405 ;
      RECT 3.295 1.725 5.02 1.895 ;
      RECT 4.72 1.35 5.02 1.725 ;
      RECT 3.51 0.925 3.68 1.725 ;
      RECT 3.175 0.595 3.68 0.925 ;
      RECT 0.115 2.37 2.665 2.54 ;
      RECT 2.495 1.8 2.665 2.37 ;
      RECT 2.495 1.47 2.785 1.8 ;
      RECT 0.115 2.54 0.445 2.83 ;
      RECT 0.115 1.95 0.855 2.37 ;
      RECT 0.685 1.28 0.855 1.95 ;
      RECT 0.115 1.11 0.855 1.28 ;
      RECT 0.115 0.61 0.445 1.11 ;
      RECT 1.185 1.95 1.63 2.2 ;
      RECT 1.46 1.78 1.63 1.95 ;
      RECT 1.46 1.45 1.9 1.78 ;
      RECT 1.46 1.2 1.63 1.45 ;
      RECT 1.24 0.94 1.63 1.2 ;
      RECT 1.24 0.77 3.005 0.94 ;
      RECT 2.835 0.425 3.005 0.77 ;
      RECT 1.24 0.42 1.63 0.77 ;
      RECT 2.835 0.255 4.02 0.425 ;
      RECT 3.85 0.425 4.02 1.225 ;
      RECT 3.85 1.225 4.15 1.555 ;
      RECT 5.19 1.62 8.595 1.63 ;
      RECT 6.765 1.3 8.595 1.62 ;
      RECT 5.19 1.63 6.935 1.79 ;
      RECT 6.11 1.79 6.44 2.7 ;
      RECT 5.11 2.48 5.44 2.7 ;
      RECT 4.195 2.065 5.44 2.48 ;
      RECT 5.19 1.79 5.44 2.065 ;
      RECT 5.19 0.95 5.36 1.62 ;
      RECT 5.18 0.62 5.36 0.95 ;
      RECT 0 -0.085 9.12 0.085 ;
      RECT 8.675 0.085 9.005 0.71 ;
      RECT 5.965 0.085 6.295 0.6 ;
      RECT 6.955 0.085 7.215 1.13 ;
      RECT 7.815 0.085 8.145 0.71 ;
      RECT 0.68 0.085 1.01 0.94 ;
      RECT 2.335 0.085 2.665 0.6 ;
      RECT 4.19 0.085 4.44 0.81 ;
      RECT 0 3.245 9.12 3.415 ;
      RECT 8.595 2.14 8.925 3.245 ;
      RECT 0.65 2.71 0.98 3.245 ;
      RECT 2.335 2.71 2.665 3.245 ;
      RECT 4.345 2.65 4.905 3.245 ;
      RECT 5.61 1.96 5.94 3.245 ;
      RECT 6.645 1.96 6.975 3.245 ;
      RECT 7.595 2.14 7.925 3.245 ;
      RECT 2.845 2.905 3.985 3.075 ;
      RECT 2.845 2.14 3.015 2.905 ;
      RECT 3.655 2.065 3.985 2.905 ;
      RECT 2.845 1.97 3.125 2.14 ;
      RECT 2.955 1.45 3.125 1.97 ;
      RECT 2.955 1.28 3.34 1.45 ;
      RECT 1.8 1.11 3.34 1.28 ;
      RECT 2.07 1.28 2.24 2.02 ;
      RECT 1.8 2.02 2.24 2.2 ;
    LAYER mcon ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
  END
END scs8ls_dlrtp_4

MACRO scs8ls_dlxbn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN GATEN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.69 1.335 2.15 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END GATEN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.79 0.35 6.13 1.1 ;
        RECT 5.96 1.1 6.13 1.82 ;
        RECT 5.765 1.82 6.13 2.98 ;
    END
    ANTENNADIFFAREA 0.5245 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.715 0.35 8.05 2.98 ;
    END
    ANTENNADIFFAREA 0.5376 ;
  END QN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.26 0.835 1.93 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.845 1.88 2.91 2.22 ;
      RECT 2.075 1.71 3.34 1.88 ;
      RECT 3.035 1.47 3.34 1.71 ;
      RECT 2.075 1.09 2.245 1.71 ;
      RECT 3.035 0.505 3.205 1.47 ;
      RECT 1.695 0.92 2.245 1.09 ;
      RECT 3.035 0.255 4.26 0.505 ;
      RECT 1.235 2.56 1.565 2.98 ;
      RECT 1.235 2.39 4.145 2.56 ;
      RECT 1.235 2.32 1.675 2.39 ;
      RECT 3.975 1.8 4.145 2.39 ;
      RECT 1.505 1.52 1.675 2.32 ;
      RECT 3.85 1.47 4.145 1.8 ;
      RECT 1.135 1.26 1.905 1.52 ;
      RECT 1.135 0.92 1.465 1.26 ;
      RECT 5.39 1.27 5.79 1.6 ;
      RECT 5.22 1.89 5.56 2.9 ;
      RECT 4.315 1.72 5.56 1.89 ;
      RECT 5.39 1.6 5.56 1.72 ;
      RECT 4.315 1.47 4.645 1.72 ;
      RECT 5.39 0.96 5.56 1.27 ;
      RECT 5.205 0.35 5.56 0.96 ;
      RECT 6.72 1.63 7.065 2.98 ;
      RECT 6.72 1.3 7.5 1.63 ;
      RECT 6.72 0.54 7.06 1.3 ;
      RECT 0.095 0.58 2.865 0.75 ;
      RECT 2.535 0.75 2.865 1.51 ;
      RECT 0.095 2.1 0.545 2.98 ;
      RECT 0.095 0.75 0.445 1.09 ;
      RECT 0.095 1.09 0.265 2.1 ;
      RECT 3.26 2.05 3.805 2.22 ;
      RECT 3.51 1.3 3.68 2.05 ;
      RECT 3.51 1.13 5.22 1.3 ;
      RECT 4.89 1.3 5.22 1.55 ;
      RECT 3.51 1.055 4.135 1.13 ;
      RECT 3.375 0.725 4.135 1.055 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 6.3 2.1 6.55 3.245 ;
      RECT 7.265 1.82 7.515 3.245 ;
      RECT 2.38 2.73 2.71 3.245 ;
      RECT 0.735 2.32 1.065 3.245 ;
      RECT 4.48 2.06 5.02 3.245 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 6.3 0.085 6.55 1.13 ;
      RECT 7.29 0.085 7.54 1.13 ;
      RECT 0.625 0.085 0.955 0.41 ;
      RECT 2.34 0.085 2.675 0.41 ;
      RECT 4.705 0.085 5.035 0.96 ;
    LAYER mcon ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
  END
END scs8ls_dlxbn_1

MACRO scs8ls_dlxbn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.225 1.82 8.555 2.98 ;
        RECT 8.325 1.13 8.495 1.82 ;
        RECT 8.245 0.35 8.495 1.13 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.13 6.115 1.8 ;
        RECT 5.885 1.8 6.59 2.07 ;
        RECT 5.885 0.85 6.505 1.13 ;
        RECT 6.245 0.355 6.505 0.85 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END Q

  PIN GATEN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.985 1.695 1.315 2.15 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END GATEN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.44 1.45 0.815 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 5.25 2.24 6.955 2.41 ;
      RECT 6.785 1.63 6.955 2.24 ;
      RECT 6.285 1.3 6.955 1.63 ;
      RECT 5.25 2.41 5.655 2.98 ;
      RECT 5.25 1.89 5.655 2.24 ;
      RECT 4.445 1.72 5.655 1.89 ;
      RECT 4.445 1.355 4.775 1.72 ;
      RECT 5.485 0.845 5.655 1.72 ;
      RECT 5.185 0.35 5.655 0.845 ;
      RECT 7.215 1.65 7.545 2.98 ;
      RECT 7.215 1.32 8.155 1.65 ;
      RECT 7.215 1.13 7.515 1.32 ;
      RECT 7.185 0.45 7.515 1.13 ;
      RECT 1.825 1.88 2.155 2.22 ;
      RECT 1.825 1.71 3.385 1.88 ;
      RECT 3.015 1.47 3.385 1.71 ;
      RECT 2.055 1.09 2.225 1.71 ;
      RECT 3.015 0.505 3.185 1.47 ;
      RECT 1.695 0.92 2.225 1.09 ;
      RECT 3.015 0.255 4.265 0.505 ;
      RECT 0.1 0.58 2.845 0.75 ;
      RECT 2.515 0.75 2.845 1.54 ;
      RECT 0.1 2.1 0.445 2.98 ;
      RECT 0.1 0.75 0.445 1.25 ;
      RECT 0.1 1.25 0.27 2.1 ;
      RECT 1.15 2.56 1.485 2.98 ;
      RECT 1.15 2.39 4.275 2.56 ;
      RECT 1.15 2.32 1.655 2.39 ;
      RECT 4.105 1.75 4.275 2.39 ;
      RECT 1.485 1.525 1.655 2.32 ;
      RECT 3.895 1.42 4.275 1.75 ;
      RECT 1.135 1.26 1.885 1.525 ;
      RECT 1.135 0.92 1.465 1.26 ;
      RECT 0 -0.085 9.12 0.085 ;
      RECT 8.675 0.085 9.005 1.13 ;
      RECT 6.675 0.085 7.005 1.13 ;
      RECT 7.745 0.085 8.075 1.13 ;
      RECT 0.625 0.085 0.955 0.41 ;
      RECT 2.285 0.085 2.64 0.41 ;
      RECT 4.63 0.085 5.015 0.845 ;
      RECT 5.825 0.085 6.075 0.68 ;
      RECT 0 3.245 9.12 3.415 ;
      RECT 8.755 1.82 9.005 3.245 ;
      RECT 5.89 2.58 6.14 3.245 ;
      RECT 6.71 2.58 7.04 3.245 ;
      RECT 7.775 1.82 8.025 3.245 ;
      RECT 2.36 2.73 2.69 3.245 ;
      RECT 4.67 2.07 5.08 3.245 ;
      RECT 0.65 2.32 0.98 3.245 ;
      RECT 3.23 2.05 3.935 2.22 ;
      RECT 3.555 1.185 3.725 2.05 ;
      RECT 3.555 1.055 5.315 1.185 ;
      RECT 4.985 1.185 5.315 1.55 ;
      RECT 3.355 1.015 5.315 1.055 ;
      RECT 3.355 0.725 4.07 1.015 ;
    LAYER mcon ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
  END
END scs8ls_dlxbn_2

MACRO scs8ls_dlxbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435 1.22 0.835 1.89 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END D

  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.18 1.335 1.55 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END GATE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.795 0.37 6.125 1.15 ;
        RECT 5.955 1.15 6.125 1.82 ;
        RECT 5.765 1.82 6.125 2.98 ;
    END
    ANTENNADIFFAREA 0.5376 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.715 0.35 8.05 2.98 ;
    END
    ANTENNADIFFAREA 0.5357 ;
  END QN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.93 2.61 2.18 2.82 ;
      RECT 1.93 2.44 4.1 2.61 ;
      RECT 1.93 2.4 2.18 2.44 ;
      RECT 3.77 2.05 4.1 2.44 ;
      RECT 3.045 1.48 3.215 2.44 ;
      RECT 3.045 1.19 3.515 1.48 ;
      RECT 1.845 1.02 3.515 1.19 ;
      RECT 1.845 0.92 2.175 1.02 ;
      RECT 1.17 1.89 1.42 2.375 ;
      RECT 1.17 1.72 2.33 1.89 ;
      RECT 1.505 1.47 2.33 1.72 ;
      RECT 1.505 1.01 1.675 1.47 ;
      RECT 1.13 0.75 1.675 1.01 ;
      RECT 1.13 0.58 3.08 0.75 ;
      RECT 2.91 0.51 3.08 0.58 ;
      RECT 1.13 0.35 1.675 0.58 ;
      RECT 2.91 0.255 4.075 0.51 ;
      RECT 0.095 2.545 1.76 2.715 ;
      RECT 1.59 2.23 1.76 2.545 ;
      RECT 1.59 2.06 2.875 2.23 ;
      RECT 2.545 1.47 2.875 2.06 ;
      RECT 0.095 2.715 0.44 2.925 ;
      RECT 0.095 2.06 0.44 2.545 ;
      RECT 0.095 0.54 0.45 1.05 ;
      RECT 0.095 1.05 0.265 2.06 ;
      RECT 5.205 1.32 5.775 1.65 ;
      RECT 5.205 2.32 5.535 2.98 ;
      RECT 4.315 1.99 5.535 2.32 ;
      RECT 5.205 1.65 5.535 1.99 ;
      RECT 5.205 1.07 5.375 1.32 ;
      RECT 5.02 0.35 5.375 1.07 ;
      RECT 6.72 1.65 7.05 2.98 ;
      RECT 6.72 1.32 7.32 1.65 ;
      RECT 6.72 0.56 7.055 1.32 ;
      RECT 3.385 1.82 3.555 2.27 ;
      RECT 3.385 1.65 5.035 1.82 ;
      RECT 4.705 1.24 5.035 1.65 ;
      RECT 3.78 0.85 3.95 1.65 ;
      RECT 3.31 0.68 3.95 0.85 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 6.295 2.1 6.545 3.245 ;
      RECT 7.27 1.82 7.52 3.245 ;
      RECT 0.64 2.885 0.97 3.245 ;
      RECT 2.38 2.78 2.71 3.245 ;
      RECT 4.49 2.545 5.035 3.245 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 6.295 0.085 6.545 1.15 ;
      RECT 7.285 0.085 7.535 1.13 ;
      RECT 0.63 0.085 0.96 1.01 ;
      RECT 2.355 0.085 2.74 0.41 ;
      RECT 4.52 0.085 4.85 1.06 ;
    LAYER mcon ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
  END
END scs8ls_dlxbp_1

MACRO scs8ls_dlxtn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.435 1.565 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END D

  PIN GATEN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.945 1.5 1.315 1.83 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END GATEN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.27 0.35 6.605 2.98 ;
    END
    ANTENNADIFFAREA 0.545 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.33 2.065 3.84 2.735 ;
      RECT 3.67 1.055 3.84 2.065 ;
      RECT 3.655 0.805 4.68 1.055 ;
      RECT 4.51 1.055 4.68 1.305 ;
      RECT 4.51 1.305 5.315 1.635 ;
      RECT 5.265 2.355 5.655 2.98 ;
      RECT 4.35 2.025 5.655 2.355 ;
      RECT 5.265 1.94 5.655 2.025 ;
      RECT 5.485 1.63 5.655 1.94 ;
      RECT 5.485 1.3 5.885 1.63 ;
      RECT 5.485 1.135 5.655 1.3 ;
      RECT 5.28 0.455 5.655 1.135 ;
      RECT 1.155 2.61 1.655 2.955 ;
      RECT 1.155 2.44 3.045 2.61 ;
      RECT 2.875 2.61 3.045 2.905 ;
      RECT 1.155 2.075 1.655 2.44 ;
      RECT 2.875 2.905 4.18 3.075 ;
      RECT 1.485 1.77 1.655 2.075 ;
      RECT 4.01 1.785 4.18 2.905 ;
      RECT 1.485 1.33 1.885 1.77 ;
      RECT 4.01 1.455 4.34 1.785 ;
      RECT 1.135 1 1.885 1.33 ;
      RECT 1.485 0.76 1.885 1 ;
      RECT 1.825 1.94 2.225 2.27 ;
      RECT 2.055 1.895 2.225 1.94 ;
      RECT 2.055 1.725 3.5 1.895 ;
      RECT 3.18 1.47 3.5 1.725 ;
      RECT 2.055 0.595 2.305 1.725 ;
      RECT 3.315 0.585 3.485 1.47 ;
      RECT 3.315 0.255 4.355 0.585 ;
      RECT 0.115 0.66 1.315 0.83 ;
      RECT 1.145 0.425 1.315 0.66 ;
      RECT 1.145 0.255 2.645 0.425 ;
      RECT 2.475 0.425 2.645 1.225 ;
      RECT 2.475 1.225 2.97 1.555 ;
      RECT 0.12 1.905 0.45 2.955 ;
      RECT 0.12 1.735 0.775 1.905 ;
      RECT 0.605 1.01 0.775 1.735 ;
      RECT 0.115 0.83 0.775 1.01 ;
      RECT 0.115 0.555 0.445 0.66 ;
      RECT 0 3.245 6.72 3.415 ;
      RECT 2.36 2.78 2.705 3.245 ;
      RECT 4.47 2.525 5.065 3.245 ;
      RECT 0.62 2.075 0.95 3.245 ;
      RECT 5.825 1.82 6.075 3.245 ;
      RECT 0 -0.085 6.72 0.085 ;
      RECT 0.625 0.085 0.955 0.49 ;
      RECT 2.815 0.085 3.145 1.055 ;
      RECT 4.85 0.085 5.1 1.135 ;
      RECT 5.84 0.085 6.09 1.13 ;
    LAYER mcon ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
  END
END scs8ls_dlxtn_1

MACRO scs8ls_dlxtn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.26 1.92 6.635 2.89 ;
        RECT 6.415 1.125 6.585 1.92 ;
        RECT 6.32 0.35 6.585 1.125 ;
    END
    ANTENNADIFFAREA 0.638 ;
  END Q

  PIN GATEN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.985 1.45 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.237 ;
  END GATEN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.3 0.455 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 5.25 2.355 5.58 2.955 ;
      RECT 4.36 2.025 5.58 2.355 ;
      RECT 5.25 1.965 5.58 2.025 ;
      RECT 5.25 1.795 5.675 1.965 ;
      RECT 5.505 1.625 5.675 1.795 ;
      RECT 5.505 1.295 6.245 1.625 ;
      RECT 5.505 1.125 5.675 1.295 ;
      RECT 5.33 0.955 5.675 1.125 ;
      RECT 5.33 0.355 5.58 0.955 ;
      RECT 1.825 1.97 2.225 2.27 ;
      RECT 1.825 1.94 3.51 1.97 ;
      RECT 2.055 1.8 3.51 1.94 ;
      RECT 3.18 1.47 3.51 1.8 ;
      RECT 2.055 0.595 2.305 1.8 ;
      RECT 3.315 0.585 3.485 1.47 ;
      RECT 3.315 0.255 4.375 0.585 ;
      RECT 1.265 2.61 1.655 2.98 ;
      RECT 1.265 2.44 3.045 2.61 ;
      RECT 2.875 2.61 3.045 2.905 ;
      RECT 1.265 2.1 1.655 2.44 ;
      RECT 2.875 2.905 4.19 3.075 ;
      RECT 1.485 1.77 1.655 2.1 ;
      RECT 4.02 1.815 4.19 2.905 ;
      RECT 1.485 1.17 1.885 1.77 ;
      RECT 4.02 1.485 4.35 1.815 ;
      RECT 1.135 0.92 1.885 1.17 ;
      RECT 1.485 0.76 1.885 0.92 ;
      RECT 3.33 2.14 3.85 2.735 ;
      RECT 3.68 1.055 3.85 2.14 ;
      RECT 3.655 0.805 4.25 1.055 ;
      RECT 4.08 1.055 4.25 1.145 ;
      RECT 4.08 1.145 5.16 1.295 ;
      RECT 4.08 1.295 5.335 1.315 ;
      RECT 4.99 1.315 5.335 1.625 ;
      RECT 0 -0.085 7.2 0.085 ;
      RECT 6.755 0.085 7.085 1.13 ;
      RECT 0.625 0.085 0.955 0.41 ;
      RECT 2.815 0.085 3.145 1.055 ;
      RECT 4.82 0.085 5.15 0.975 ;
      RECT 5.845 0.085 6.14 1.125 ;
      RECT 0 3.245 7.2 3.415 ;
      RECT 6.835 1.82 7.085 3.245 ;
      RECT 2.36 2.78 2.705 3.245 ;
      RECT 4.36 2.625 5.08 3.245 ;
      RECT 0.765 2.29 1.095 3.245 ;
      RECT 5.845 1.82 6.06 3.245 ;
      RECT 0.115 0.58 1.315 0.75 ;
      RECT 1.145 0.425 1.315 0.58 ;
      RECT 1.145 0.255 2.645 0.425 ;
      RECT 2.475 0.425 2.645 1.3 ;
      RECT 2.475 1.3 2.97 1.63 ;
      RECT 0.265 2.12 0.595 2.98 ;
      RECT 0.265 1.95 0.795 2.12 ;
      RECT 0.625 1.13 0.795 1.95 ;
      RECT 0.115 0.75 0.795 1.13 ;
    LAYER mcon ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
  END
END scs8ls_dlxtn_2

MACRO scs8ls_clkbuf_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.095 1.78 ;
    END
    ANTENNAGATEAREA 0.462 ;
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.71 1.18 5.155 1.69 ;
        RECT 1.615 1.69 5.155 1.86 ;
        RECT 4.71 1.02 4.88 1.18 ;
        RECT 1.615 1.86 1.88 2.98 ;
        RECT 2.585 1.86 2.845 2.98 ;
        RECT 3.415 1.86 3.68 2.98 ;
        RECT 4.385 1.86 4.645 2.98 ;
        RECT 1.615 0.85 4.88 1.02 ;
        RECT 1.615 0.35 1.945 0.85 ;
        RECT 2.615 0.35 2.865 0.85 ;
        RECT 3.555 0.35 3.725 0.85 ;
        RECT 4.485 0.35 4.655 0.85 ;
    END
    ANTENNADIFFAREA 1.8417 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.275 1.19 4.515 1.52 ;
      RECT 0.615 2.12 0.945 2.98 ;
      RECT 0.615 1.95 1.445 2.12 ;
      RECT 1.275 1.52 1.445 1.95 ;
      RECT 1.275 1.15 1.445 1.19 ;
      RECT 0.615 0.98 1.445 1.15 ;
      RECT 0.615 0.35 0.945 0.98 ;
      RECT 0 3.245 5.28 3.415 ;
      RECT 4.83 2.03 5.16 3.245 ;
      RECT 1.115 2.29 1.445 3.245 ;
      RECT 0.115 1.95 0.445 3.245 ;
      RECT 2.065 2.03 2.395 3.245 ;
      RECT 3.045 2.03 3.215 3.245 ;
      RECT 3.865 2.03 4.195 3.245 ;
      RECT 0 -0.085 5.28 0.085 ;
      RECT 4.835 0.085 5.165 0.68 ;
      RECT 0.115 0.085 0.445 0.81 ;
      RECT 1.115 0.085 1.445 0.81 ;
      RECT 2.115 0.085 2.445 0.68 ;
      RECT 3.045 0.085 3.375 0.68 ;
      RECT 3.905 0.085 4.305 0.68 ;
    LAYER mcon ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_clkbuf_8

MACRO scs8ls_clkdlyinv3sd1_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.53 0.755 2.795 1.815 ;
        RECT 2.435 1.815 2.795 3.06 ;
        RECT 2.435 0.355 2.795 0.755 ;
    END
    ANTENNADIFFAREA 0.4249 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.19 0.73 1.86 ;
    END
    ANTENNAGATEAREA 0.231 ;
  END A

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.88 0.085 ;
      RECT 0.585 0.085 0.915 0.65 ;
      RECT 1.935 0.085 2.265 0.75 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 0.575 2.38 0.905 3.245 ;
      RECT 1.935 1.9 2.265 3.245 ;
      RECT 1.415 2.65 1.745 2.9 ;
      RECT 1.475 1.625 1.745 2.65 ;
      RECT 1.475 1.295 2.36 1.625 ;
      RECT 1.475 0.305 1.72 1.295 ;
      RECT 0.095 2.205 0.4 2.725 ;
      RECT 0.095 2.03 1.305 2.205 ;
      RECT 0.975 1.02 1.305 2.03 ;
      RECT 0.095 0.82 1.305 1.02 ;
      RECT 0.095 0.305 0.41 0.82 ;
    LAYER mcon ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_clkdlyinv3sd1_1

MACRO scs8ls_clkdlyinv3sd2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.53 0.755 2.795 1.815 ;
        RECT 2.435 1.815 2.795 3.06 ;
        RECT 2.435 0.355 2.795 0.755 ;
    END
    ANTENNADIFFAREA 0.4249 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.19 0.73 1.86 ;
    END
    ANTENNAGATEAREA 0.231 ;
  END A

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.88 0.085 ;
      RECT 0.585 0.085 0.915 0.65 ;
      RECT 1.935 0.085 2.265 0.75 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 0.575 2.38 0.905 3.245 ;
      RECT 1.935 1.9 2.265 3.245 ;
      RECT 1.415 2.65 1.745 2.9 ;
      RECT 1.475 1.625 1.745 2.65 ;
      RECT 1.475 1.295 2.36 1.625 ;
      RECT 1.475 0.305 1.72 1.295 ;
      RECT 0.095 2.205 0.4 2.725 ;
      RECT 0.095 2.03 1.305 2.205 ;
      RECT 0.975 1.02 1.305 2.03 ;
      RECT 0.095 0.82 1.305 1.02 ;
      RECT 0.095 0.305 0.41 0.82 ;
    LAYER mcon ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_clkdlyinv3sd2_1

MACRO scs8ls_clkdlyinv3sd3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.53 0.755 2.795 1.815 ;
        RECT 2.435 1.815 2.795 3.06 ;
        RECT 2.435 0.355 2.795 0.755 ;
    END
    ANTENNADIFFAREA 0.4249 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.19 0.73 1.86 ;
    END
    ANTENNAGATEAREA 0.231 ;
  END A

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 2.88 0.085 ;
      RECT 0.585 0.085 0.915 0.65 ;
      RECT 1.935 0.085 2.265 0.75 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 0.575 2.38 0.905 3.245 ;
      RECT 1.935 1.9 2.265 3.245 ;
      RECT 1.415 2.65 1.745 2.9 ;
      RECT 1.475 1.625 1.745 2.65 ;
      RECT 1.475 1.295 2.36 1.625 ;
      RECT 1.475 0.305 1.72 1.295 ;
      RECT 0.095 2.205 0.4 2.725 ;
      RECT 0.095 2.03 1.305 2.205 ;
      RECT 0.975 1.02 1.305 2.03 ;
      RECT 0.095 0.82 1.305 1.02 ;
      RECT 0.095 0.305 0.41 0.82 ;
    LAYER mcon ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_clkdlyinv3sd3_1

MACRO scs8ls_clkdlyinv5sd1_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 0.755 5.19 1.9 ;
        RECT 4.83 1.9 5.19 3.06 ;
        RECT 4.83 0.355 5.19 0.755 ;
    END
    ANTENNADIFFAREA 0.4249 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.19 0.73 1.86 ;
    END
    ANTENNAGATEAREA 0.231 ;
  END A

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.415 1.73 3.655 2.98 ;
      RECT 3.415 1.56 4.755 1.73 ;
      RECT 4.53 1.05 4.755 1.56 ;
      RECT 3.37 0.925 4.755 1.05 ;
      RECT 3.37 0.88 4.7 0.925 ;
      RECT 3.37 0.4 3.7 0.88 ;
      RECT 2.8 1.39 2.97 2.98 ;
      RECT 2.8 1.22 4.005 1.39 ;
      RECT 2.8 0.415 2.97 1.22 ;
      RECT 0 3.245 5.28 3.415 ;
      RECT 0.575 2.38 0.905 3.245 ;
      RECT 1.915 1.94 2.265 3.245 ;
      RECT 4.33 1.9 4.66 3.245 ;
      RECT 1.415 2.65 1.745 2.9 ;
      RECT 1.475 1.47 1.745 2.65 ;
      RECT 1.475 1.14 2.51 1.47 ;
      RECT 1.475 0.305 1.72 1.14 ;
      RECT 0 -0.085 5.28 0.085 ;
      RECT 0.585 0.085 0.915 0.65 ;
      RECT 1.915 0.085 2.265 0.745 ;
      RECT 4.33 0.085 4.66 0.67 ;
      RECT 0.095 2.205 0.4 2.725 ;
      RECT 0.095 2.03 1.305 2.205 ;
      RECT 0.975 1.02 1.305 2.03 ;
      RECT 0.095 0.82 1.305 1.02 ;
      RECT 0.095 0.305 0.41 0.82 ;
    LAYER mcon ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
  END
END scs8ls_clkdlyinv5sd1_1

MACRO scs8ls_clkdlyinv5sd2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 0.755 5.19 1.9 ;
        RECT 4.83 1.9 5.19 3.06 ;
        RECT 4.83 0.355 5.19 0.755 ;
    END
    ANTENNADIFFAREA 0.4249 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.19 0.73 1.86 ;
    END
    ANTENNAGATEAREA 0.231 ;
  END A

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.415 1.73 3.655 2.98 ;
      RECT 3.415 1.56 4.755 1.73 ;
      RECT 4.53 1.05 4.755 1.56 ;
      RECT 3.37 0.925 4.755 1.05 ;
      RECT 3.37 0.88 4.7 0.925 ;
      RECT 3.37 0.4 3.7 0.88 ;
      RECT 2.8 1.39 2.97 2.98 ;
      RECT 2.8 1.22 4.005 1.39 ;
      RECT 2.8 0.415 2.97 1.22 ;
      RECT 0 3.245 5.28 3.415 ;
      RECT 0.575 2.38 0.905 3.245 ;
      RECT 1.915 1.94 2.265 3.245 ;
      RECT 4.33 1.9 4.66 3.245 ;
      RECT 1.415 2.65 1.745 2.9 ;
      RECT 1.475 1.47 1.745 2.65 ;
      RECT 1.475 1.14 2.51 1.47 ;
      RECT 1.475 0.305 1.72 1.14 ;
      RECT 0 -0.085 5.28 0.085 ;
      RECT 0.585 0.085 0.915 0.65 ;
      RECT 1.915 0.085 2.265 0.745 ;
      RECT 4.33 0.085 4.66 0.67 ;
      RECT 0.095 2.205 0.4 2.725 ;
      RECT 0.095 2.03 1.305 2.205 ;
      RECT 0.975 1.02 1.305 2.03 ;
      RECT 0.095 0.82 1.305 1.02 ;
      RECT 0.095 0.305 0.41 0.82 ;
    LAYER mcon ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
  END
END scs8ls_clkdlyinv5sd2_1

MACRO scs8ls_clkdlyinv5sd3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 0.755 5.19 1.9 ;
        RECT 4.83 1.9 5.19 3.06 ;
        RECT 4.83 0.355 5.19 0.755 ;
    END
    ANTENNADIFFAREA 0.4249 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.19 0.73 1.86 ;
    END
    ANTENNAGATEAREA 0.231 ;
  END A

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.415 1.73 3.655 2.98 ;
      RECT 3.415 1.56 4.755 1.73 ;
      RECT 4.53 1.05 4.755 1.56 ;
      RECT 3.37 0.925 4.755 1.05 ;
      RECT 3.37 0.88 4.7 0.925 ;
      RECT 3.37 0.4 3.7 0.88 ;
      RECT 2.8 1.39 2.97 2.98 ;
      RECT 2.8 1.22 4.005 1.39 ;
      RECT 2.8 0.415 2.97 1.22 ;
      RECT 0 3.245 5.28 3.415 ;
      RECT 0.575 2.38 0.905 3.245 ;
      RECT 1.915 1.94 2.265 3.245 ;
      RECT 4.33 1.9 4.66 3.245 ;
      RECT 1.415 2.65 1.745 2.9 ;
      RECT 1.475 1.47 1.745 2.65 ;
      RECT 1.475 1.14 2.51 1.47 ;
      RECT 1.475 0.305 1.72 1.14 ;
      RECT 0 -0.085 5.28 0.085 ;
      RECT 0.585 0.085 0.915 0.65 ;
      RECT 1.915 0.085 2.265 0.745 ;
      RECT 4.33 0.085 4.66 0.67 ;
      RECT 0.095 2.205 0.4 2.725 ;
      RECT 0.095 2.03 1.305 2.205 ;
      RECT 0.975 1.02 1.305 2.03 ;
      RECT 0.095 0.82 1.305 1.02 ;
      RECT 0.095 0.305 0.41 0.82 ;
    LAYER mcon ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
  END
END scs8ls_clkdlyinv5sd3_1

MACRO scs8ls_clkinv_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615 0.35 1.325 0.68 ;
        RECT 1.085 0.68 1.325 2.1 ;
        RECT 0.555 2.1 1.325 2.43 ;
        RECT 0.555 2.43 0.835 2.955 ;
    END
    ANTENNADIFFAREA 0.47735 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.755 1.78 ;
        RECT 0.425 1.78 0.755 1.93 ;
        RECT 0.425 0.92 0.755 1.18 ;
    END
    ANTENNAGATEAREA 0.315 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 1.44 0.085 ;
      RECT 0.115 0.085 0.445 0.75 ;
      RECT 0 3.245 1.44 3.415 ;
      RECT 1.005 2.6 1.335 3.245 ;
      RECT 0.105 2.1 0.355 3.245 ;
    LAYER mcon ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_clkinv_1

MACRO scs8ls_clkinv_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 11.52 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.575 1.92 10.935 2.15 ;
    END
    ANTENNADIFFAREA 5.04 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.985 1.18 10.935 1.41 ;
    END
    ANTENNAGATEAREA 5.04 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.52 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.52 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.705 1.95 10.875 2.12 ;
      RECT 10.625 1.21 10.795 1.38 ;
      RECT 10.265 1.21 10.435 1.38 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.905 1.21 10.075 1.38 ;
      RECT 9.805 1.95 9.975 2.12 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.545 1.21 9.715 1.38 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 9.185 1.21 9.355 1.38 ;
      RECT 8.905 1.95 9.075 2.12 ;
      RECT 8.825 1.21 8.995 1.38 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.465 1.21 8.635 1.38 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 8.105 1.21 8.275 1.38 ;
      RECT 8.005 1.95 8.175 2.12 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.745 1.21 7.915 1.38 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.075 1.95 7.245 2.12 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.625 1.21 6.795 1.38 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 6.095 1.95 6.265 2.12 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.675 1.21 5.845 1.38 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 5.145 1.95 5.315 2.12 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.835 1.21 5.005 1.38 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.245 1.95 4.415 2.12 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.845 1.21 4.015 1.38 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.375 1.95 3.545 2.12 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.915 1.21 3.085 1.38 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.445 1.95 2.615 2.12 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.945 1.21 2.115 1.38 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.545 1.95 1.715 2.12 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.045 1.21 1.215 1.38 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 1.95 0.805 2.12 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
    LAYER li1 ;
      RECT 5.065 2.01 5.395 2.98 ;
      RECT 5.065 1.85 5.425 2.01 ;
      RECT 5.255 0.775 5.425 1.85 ;
      RECT 5.255 0.38 5.525 0.775 ;
      RECT 5.595 1.15 5.925 1.65 ;
      RECT 0.115 0.085 0.445 0.84 ;
      RECT 0 -0.085 11.52 0.085 ;
      RECT 0.975 0.085 1.26 0.84 ;
      RECT 1.885 0.085 2.165 0.84 ;
      RECT 2.845 0.085 3.095 0.84 ;
      RECT 3.765 0.085 4.095 0.84 ;
      RECT 4.765 0.085 5.085 0.84 ;
      RECT 5.695 0.085 5.98 0.84 ;
      RECT 6.555 0.085 6.875 0.84 ;
      RECT 7.485 0.085 9.825 0.71 ;
      RECT 7.045 0.38 7.29 2.98 ;
      RECT 6.545 1.15 6.875 1.65 ;
      RECT 4.755 1.15 5.085 1.65 ;
      RECT 8.005 1.82 8.175 2.98 ;
      RECT 4.165 1.9 4.495 2.98 ;
      RECT 4.165 1.85 4.525 1.9 ;
      RECT 4.265 0.38 4.525 1.85 ;
      RECT 7.525 1.15 10.915 1.65 ;
      RECT 6.015 1.82 6.33 2.98 ;
      RECT 6.095 1.76 6.33 1.82 ;
      RECT 6.095 1.01 6.34 1.76 ;
      RECT 6.16 0.785 6.34 1.01 ;
      RECT 6.16 0.38 6.385 0.785 ;
      RECT 3.765 1.15 4.095 1.65 ;
      RECT 8.905 1.82 9.075 2.98 ;
      RECT 9.805 1.82 9.975 2.98 ;
      RECT 10.705 1.82 10.875 2.98 ;
      RECT 3.335 0.775 3.595 2.98 ;
      RECT 3.3 0.38 3.595 0.775 ;
      RECT 2.835 1.15 3.165 1.65 ;
      RECT 2.365 1.885 2.695 2.98 ;
      RECT 2.365 0.775 2.665 1.885 ;
      RECT 2.35 0.38 2.665 0.775 ;
      RECT 1.865 1.15 2.195 1.65 ;
      RECT 1.465 1.885 1.795 2.98 ;
      RECT 1.465 0.775 1.695 1.885 ;
      RECT 1.44 0.38 1.7 0.775 ;
      RECT 0.975 1.15 1.295 1.65 ;
      RECT 0.625 1.82 0.815 2.98 ;
      RECT 0.625 0.775 0.805 1.82 ;
      RECT 0.615 0.38 0.805 0.775 ;
      RECT 0 3.245 11.52 3.415 ;
      RECT 0.115 1.9 0.445 3.245 ;
      RECT 1.015 1.82 1.265 3.245 ;
      RECT 1.995 1.82 2.165 3.245 ;
      RECT 2.895 1.82 3.065 3.245 ;
      RECT 3.795 1.82 3.965 3.245 ;
      RECT 4.695 1.82 4.865 3.245 ;
      RECT 5.595 1.82 5.845 3.245 ;
      RECT 6.51 1.82 6.795 3.245 ;
      RECT 7.475 1.82 7.805 3.245 ;
      RECT 8.375 1.82 8.625 3.245 ;
      RECT 9.275 1.82 9.605 3.245 ;
      RECT 10.175 1.82 10.505 3.245 ;
      RECT 11.075 1.82 11.405 3.245 ;
  END
END scs8ls_clkinv_16

MACRO scs8ls_clkinv_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.63 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.18 1.795 1.95 ;
        RECT 0.12 1.95 1.795 2.12 ;
        RECT 0.615 1.01 1.795 1.18 ;
        RECT 0.12 2.12 0.45 2.98 ;
        RECT 1.02 2.12 1.35 2.98 ;
        RECT 0.615 0.51 1.305 1.01 ;
    END
    ANTENNADIFFAREA 0.994 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 1.92 3.415 ;
      RECT 1.55 2.29 1.8 3.245 ;
      RECT 0.65 2.29 0.82 3.245 ;
      RECT 0 -0.085 1.92 0.085 ;
      RECT 1.475 0.085 1.805 0.84 ;
      RECT 0.115 0.085 0.445 0.84 ;
    LAYER mcon ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_clkinv_2

MACRO scs8ls_clkinv_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.35 2.755 1.78 ;
    END
    ANTENNAGATEAREA 1.26 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.18 3.235 1.95 ;
        RECT 0.265 1.95 3.235 2.12 ;
        RECT 0.265 1.01 3.235 1.18 ;
        RECT 0.565 2.12 0.895 2.98 ;
        RECT 1.465 2.12 1.795 2.98 ;
        RECT 2.415 2.12 2.745 2.98 ;
        RECT 0.265 1.18 0.435 1.95 ;
        RECT 0.99 0.455 1.745 1.01 ;
        RECT 2.415 0.38 2.745 1.01 ;
    END
    ANTENNADIFFAREA 1.4322 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.915 2.29 3.245 3.245 ;
      RECT 0.115 2.29 0.365 3.245 ;
      RECT 1.095 2.29 1.265 3.245 ;
      RECT 1.995 2.29 2.245 3.245 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.915 0.085 3.245 0.84 ;
      RECT 0.115 0.085 0.82 0.71 ;
      RECT 1.915 0.085 2.245 0.84 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_clkinv_4

MACRO scs8ls_clkinv_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.18 6.115 1.95 ;
        RECT 0.285 1.95 6.115 2.12 ;
        RECT 0.285 1.01 6.115 1.18 ;
        RECT 0.59 2.12 0.92 2.98 ;
        RECT 1.54 2.12 1.87 2.98 ;
        RECT 2.49 2.12 2.82 2.98 ;
        RECT 3.44 2.12 3.77 2.98 ;
        RECT 4.39 2.12 4.72 2.98 ;
        RECT 5.34 2.12 5.67 2.98 ;
        RECT 0.285 1.18 0.455 1.95 ;
        RECT 0.615 0.46 2.625 1.01 ;
        RECT 3.295 0.445 3.625 1.01 ;
        RECT 4.295 0.445 4.625 1.01 ;
        RECT 5.295 0.445 5.625 1.01 ;
    END
    ANTENNADIFFAREA 3.2424 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625 1.35 5.715 1.78 ;
    END
    ANTENNAGATEAREA 2.52 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 6.24 0.085 ;
      RECT 5.795 0.085 6.125 0.775 ;
      RECT 0.115 0.085 0.445 0.775 ;
      RECT 2.795 0.085 3.125 0.775 ;
      RECT 3.795 0.085 4.125 0.775 ;
      RECT 4.795 0.085 5.125 0.775 ;
      RECT 0 3.245 6.24 3.415 ;
      RECT 5.87 2.29 6.12 3.245 ;
      RECT 0.115 2.29 0.39 3.245 ;
      RECT 1.12 2.29 1.37 3.245 ;
      RECT 2.07 2.29 2.32 3.245 ;
      RECT 3.02 2.29 3.27 3.245 ;
      RECT 3.97 2.29 4.22 3.245 ;
      RECT 4.92 2.29 5.17 3.245 ;
    LAYER mcon ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_clkinv_8

MACRO scs8ls_conb_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.845 0.395 2.335 ;
        RECT 0.085 0.255 0.615 0.845 ;
    END
    ANTENNAPARTIALMETALSIDEAREA 0.182 LAYER li1 ;
  END HI

  PIN LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055 0.995 1.355 2.485 ;
        RECT 0.825 2.485 1.355 3.075 ;
    END
    ANTENNAPARTIALMETALSIDEAREA 0.182 LAYER li1 ;
  END LO

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.825 0.085 1.155 0.825 ;
      RECT 0 -0.085 1.44 0.085 ;
      RECT 0 3.245 1.44 3.415 ;
      RECT 0.285 2.505 0.615 3.245 ;
    LAYER mcon ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_conb_1

MACRO scs8ls_decap_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.605 0.715 0.855 1.585 ;
      RECT 0.24 0.085 0.855 0.715 ;
      RECT 0 -0.085 1.92 0.085 ;
      RECT 1.425 0.085 1.68 0.715 ;
      RECT 0 3.245 1.92 3.415 ;
      RECT 0.24 2.67 0.49 3.245 ;
      RECT 1.065 2.67 1.68 3.245 ;
      RECT 1.065 1.25 1.315 2.67 ;
    LAYER mcon ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_decap_4

MACRO scs8ls_decap_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 3.05 2.295 3.3 3.245 ;
      RECT 0.565 2.285 0.815 3.245 ;
      RECT 1.46 1.25 2.395 3.245 ;
      RECT 0.8 0.81 1.13 1.585 ;
      RECT 0.565 0.085 1.13 0.81 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 1.765 0.085 2.095 0.805 ;
      RECT 2.67 0.085 3.29 0.81 ;
      RECT 2.67 0.81 3.075 1.585 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
  END
END scs8ls_decap_8

MACRO scs8ls_dfbbn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.575 1.82 11.925 2.98 ;
        RECT 11.755 1.15 11.925 1.82 ;
        RECT 11.555 0.405 11.925 1.15 ;
    END
    ANTENNADIFFAREA 0.5134 ;
  END QN

  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.3 0.495 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLKN

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.685 1.35 11.015 1.78 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END RESETB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925 1.18 2.755 1.51 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.005 0.35 13.34 2.98 ;
    END
    ANTENNADIFFAREA 0.519 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.44 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.44 3.575 ;
    END
  END vpwr

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.375 1.965 9.025 2.105 ;
        RECT 5.375 2.105 5.665 2.15 ;
        RECT 8.735 2.105 9.025 2.15 ;
        RECT 5.375 1.92 5.665 1.965 ;
        RECT 8.735 1.92 9.025 1.965 ;
    END
    ANTENNAGATEAREA 0.4695 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.541 LAYER met1 ;
  END SETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.795 1.95 8.965 2.12 ;
      RECT 6.875 1.21 7.045 1.38 ;
      RECT 5.435 1.95 5.605 2.12 ;
      RECT 3.035 1.21 3.205 1.38 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
    LAYER met1 ;
      RECT 2.975 1.365 3.265 1.41 ;
      RECT 2.975 1.225 7.105 1.365 ;
      RECT 6.815 1.365 7.105 1.41 ;
      RECT 2.975 1.18 3.265 1.225 ;
      RECT 6.815 1.18 7.105 1.225 ;
    LAYER li1 ;
      RECT 5.435 1.96 5.635 2.15 ;
      RECT 5.435 1.675 5.85 1.96 ;
      RECT 9.065 0.425 9.315 0.765 ;
      RECT 9.065 0.255 10.36 0.425 ;
      RECT 10.345 1.95 10.85 2.12 ;
      RECT 8.375 0.935 10.89 1.105 ;
      RECT 10.345 1.105 10.515 1.95 ;
      RECT 9.3 1.105 9.63 1.56 ;
      RECT 8.375 0.51 8.545 0.935 ;
      RECT 6.315 0.34 8.545 0.51 ;
      RECT 6.315 0.51 6.485 1.335 ;
      RECT 4.985 1.335 6.485 1.505 ;
      RECT 4.985 1.505 5.265 1.665 ;
      RECT 4.315 0.425 4.645 0.825 ;
      RECT 4.315 0.255 5.645 0.425 ;
      RECT 5.315 0.425 5.645 1.035 ;
      RECT 0.105 2.12 0.435 2.98 ;
      RECT 0.105 1.95 0.835 2.12 ;
      RECT 0.665 1.63 0.835 1.95 ;
      RECT 0.665 1.3 1.075 1.63 ;
      RECT 0.665 1.13 0.835 1.3 ;
      RECT 0.115 0.96 0.835 1.13 ;
      RECT 0.115 0.35 0.365 0.96 ;
      RECT 1.005 2.905 2.125 3.075 ;
      RECT 1.955 1.855 2.125 2.905 ;
      RECT 1.955 1.685 3.24 1.855 ;
      RECT 2.975 1.855 3.24 2.355 ;
      RECT 2.975 1.455 3.24 1.685 ;
      RECT 2.975 1.125 3.465 1.455 ;
      RECT 1.005 1.82 1.415 2.905 ;
      RECT 1.245 1.13 1.415 1.82 ;
      RECT 1.055 0.35 1.415 1.13 ;
      RECT 2.635 2.905 4.53 3.075 ;
      RECT 4.2 2.49 4.53 2.905 ;
      RECT 2.635 2.355 2.805 2.905 ;
      RECT 4.2 2.32 6.45 2.49 ;
      RECT 2.37 2.025 2.805 2.355 ;
      RECT 5.57 2.49 5.82 2.98 ;
      RECT 4.2 2.305 4.815 2.32 ;
      RECT 6.12 1.675 6.45 2.32 ;
      RECT 4.645 1.165 4.815 2.305 ;
      RECT 4.645 0.995 5.145 1.165 ;
      RECT 4.815 0.715 5.145 0.995 ;
      RECT 8.39 2.29 9.4 2.46 ;
      RECT 9.23 2.12 9.4 2.29 ;
      RECT 8.39 1.9 8.56 2.29 ;
      RECT 9.23 1.95 10.17 2.12 ;
      RECT 7.245 1.73 8.56 1.9 ;
      RECT 9.84 1.42 10.17 1.95 ;
      RECT 7.245 1.9 7.415 2.1 ;
      RECT 8.035 1.01 8.205 1.73 ;
      RECT 6.86 2.1 7.415 2.98 ;
      RECT 6.72 0.68 8.205 1.01 ;
      RECT 11.215 1.32 11.585 1.65 ;
      RECT 9.99 2.29 11.385 2.46 ;
      RECT 11.215 1.65 11.385 2.29 ;
      RECT 11.215 0.765 11.385 1.32 ;
      RECT 9.495 0.595 11.385 0.765 ;
      RECT 8.5 2.8 8.83 2.98 ;
      RECT 7.89 2.63 10.32 2.8 ;
      RECT 9.99 2.8 10.32 2.98 ;
      RECT 9.99 2.46 10.32 2.63 ;
      RECT 7.89 2.07 8.22 2.63 ;
      RECT 8.73 1.275 9.06 2.12 ;
      RECT 3.09 2.565 3.58 2.735 ;
      RECT 3.41 1.795 3.58 2.565 ;
      RECT 3.41 1.625 4.135 1.795 ;
      RECT 3.635 1.395 4.135 1.625 ;
      RECT 3.635 0.955 3.805 1.395 ;
      RECT 2.95 0.785 3.805 0.955 ;
      RECT 2.95 0.595 3.28 0.785 ;
      RECT 1.585 0.84 2.75 1.01 ;
      RECT 2.58 0.425 2.75 0.84 ;
      RECT 2.58 0.255 4.145 0.425 ;
      RECT 3.46 0.425 4.145 0.615 ;
      RECT 3.975 0.615 4.145 0.995 ;
      RECT 3.975 0.995 4.475 1.165 ;
      RECT 4.305 1.165 4.475 1.965 ;
      RECT 3.75 1.965 4.475 2.135 ;
      RECT 3.75 2.135 4 2.735 ;
      RECT 1.585 2.405 1.785 2.735 ;
      RECT 1.585 1.01 1.755 2.405 ;
      RECT 1.585 0.575 1.865 0.84 ;
      RECT 6.71 1.56 7.075 1.93 ;
      RECT 6.71 1.18 7.865 1.56 ;
      RECT 12.11 1.585 12.36 2.91 ;
      RECT 12.11 1.255 12.835 1.585 ;
      RECT 12.11 0.35 12.36 1.255 ;
      RECT 0 -0.085 13.44 0.085 ;
      RECT 12.58 0.085 12.83 0.81 ;
      RECT 0.545 0.085 0.875 0.79 ;
      RECT 2.045 0.085 2.41 0.67 ;
      RECT 5.815 0.085 6.145 1.035 ;
      RECT 8.715 0.085 8.885 0.765 ;
      RECT 11.055 0.085 11.385 0.425 ;
      RECT 0 3.245 13.44 3.415 ;
      RECT 12.555 1.82 12.805 3.245 ;
      RECT 7.905 2.97 8.27 3.245 ;
      RECT 9.035 2.97 9.365 3.245 ;
      RECT 5.04 2.66 5.37 3.245 ;
      RECT 6.02 2.66 6.35 3.245 ;
      RECT 11.045 2.63 11.375 3.245 ;
      RECT 2.295 2.525 2.465 3.245 ;
      RECT 0.635 2.29 0.805 3.245 ;
  END
END scs8ls_dfbbn_1

MACRO scs8ls_dfbbn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 14.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.515 1.94 13.845 2.98 ;
        RECT 13.515 1.77 14.035 1.94 ;
        RECT 13.865 1.1 14.035 1.77 ;
        RECT 13.54 0.85 14.035 1.1 ;
        RECT 13.54 0.35 13.8 0.85 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.63 0.44 11.985 1.18 ;
        RECT 11.815 1.18 11.985 1.85 ;
        RECT 11.645 1.85 11.985 2.02 ;
        RECT 11.645 2.02 11.815 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END QN

  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.3 0.495 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLKN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955 1.18 2.755 1.51 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END D

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.715 1.35 11.115 1.78 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END RESETB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.4 3.575 ;
    END
  END vpwr

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.375 1.965 9.025 2.105 ;
        RECT 5.375 2.105 5.665 2.15 ;
        RECT 8.735 2.105 9.025 2.15 ;
        RECT 5.375 1.92 5.665 1.965 ;
        RECT 8.735 1.92 9.025 1.965 ;
    END
    ANTENNAGATEAREA 0.4695 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.541 LAYER met1 ;
  END SETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 1.95 5.605 2.12 ;
      RECT 8.795 1.95 8.965 2.12 ;
      RECT 6.875 1.21 7.045 1.38 ;
      RECT 3.035 1.21 3.205 1.38 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.115 -0.085 13.285 0.085 ;
    LAYER met1 ;
      RECT 2.975 1.365 3.265 1.41 ;
      RECT 2.975 1.225 7.105 1.365 ;
      RECT 6.815 1.365 7.105 1.41 ;
      RECT 2.975 1.18 3.265 1.225 ;
      RECT 6.815 1.18 7.105 1.225 ;
    LAYER li1 ;
      RECT 5.415 1.63 5.745 2.15 ;
      RECT 4.395 0.435 4.565 0.955 ;
      RECT 4.395 0.265 5.575 0.435 ;
      RECT 5.245 0.435 5.575 1.025 ;
      RECT 9.135 0.425 9.385 0.84 ;
      RECT 9.135 0.255 10.44 0.425 ;
      RECT 10.11 0.425 10.44 0.5 ;
      RECT 2.635 2.905 4.605 3.075 ;
      RECT 4.185 2.49 4.605 2.905 ;
      RECT 2.635 2.355 2.805 2.905 ;
      RECT 4.185 2.32 6.38 2.49 ;
      RECT 2.365 2.025 2.805 2.355 ;
      RECT 5.565 2.49 5.895 2.98 ;
      RECT 4.185 2.305 4.775 2.32 ;
      RECT 6.05 1.63 6.38 2.32 ;
      RECT 4.605 1.295 4.775 2.305 ;
      RECT 4.605 1.125 4.905 1.295 ;
      RECT 4.735 1.12 4.905 1.125 ;
      RECT 4.735 0.605 5.075 1.12 ;
      RECT 11.29 1.35 11.645 1.68 ;
      RECT 10.06 2.29 11.46 2.46 ;
      RECT 11.29 1.68 11.46 2.29 ;
      RECT 11.29 0.84 11.46 1.35 ;
      RECT 9.605 0.67 11.46 0.84 ;
      RECT 8.57 2.8 8.9 2.98 ;
      RECT 7.925 2.63 10.39 2.8 ;
      RECT 10.06 2.8 10.39 2.98 ;
      RECT 10.06 2.46 10.39 2.63 ;
      RECT 7.925 2.06 8.255 2.63 ;
      RECT 9.605 0.595 9.935 0.67 ;
      RECT 6.965 2.1 7.455 2.98 ;
      RECT 7.285 1.89 7.455 2.1 ;
      RECT 7.285 1.72 8.595 1.89 ;
      RECT 8.425 1.89 8.595 2.29 ;
      RECT 8.105 1.01 8.275 1.72 ;
      RECT 8.425 2.29 9.89 2.46 ;
      RECT 6.65 0.68 8.275 1.01 ;
      RECT 9.72 1.89 9.89 2.29 ;
      RECT 9.72 1.72 10.205 1.89 ;
      RECT 9.91 1.47 10.205 1.72 ;
      RECT 10.375 1.95 10.92 2.12 ;
      RECT 8.445 1.01 10.99 1.18 ;
      RECT 10.375 1.18 10.545 1.95 ;
      RECT 9.37 1.18 9.7 1.55 ;
      RECT 8.445 0.51 8.615 1.01 ;
      RECT 6.245 0.34 8.615 0.51 ;
      RECT 6.245 0.51 6.415 1.29 ;
      RECT 5.075 1.29 6.415 1.46 ;
      RECT 5.075 1.46 5.245 1.61 ;
      RECT 4.945 1.61 5.245 1.94 ;
      RECT 6.785 1.41 7.115 1.91 ;
      RECT 6.785 1.18 7.935 1.41 ;
      RECT 7.685 1.41 7.935 1.55 ;
      RECT 0.105 2.12 0.435 2.98 ;
      RECT 0.105 1.95 0.835 2.12 ;
      RECT 0.665 1.63 0.835 1.95 ;
      RECT 0.665 1.3 1.105 1.63 ;
      RECT 0.665 1.13 0.835 1.3 ;
      RECT 0.115 0.96 0.835 1.13 ;
      RECT 0.115 0.35 0.365 0.96 ;
      RECT 3.085 2.565 3.57 2.735 ;
      RECT 3.4 1.795 3.57 2.565 ;
      RECT 3.4 1.625 4.095 1.795 ;
      RECT 3.715 1.465 4.095 1.625 ;
      RECT 3.715 0.955 3.885 1.465 ;
      RECT 2.98 0.785 3.885 0.955 ;
      RECT 2.98 0.595 3.31 0.785 ;
      RECT 3.74 2.135 3.99 2.735 ;
      RECT 3.74 1.965 4.435 2.135 ;
      RECT 4.265 1.295 4.435 1.965 ;
      RECT 4.055 1.125 4.435 1.295 ;
      RECT 4.055 0.615 4.225 1.125 ;
      RECT 3.49 0.425 4.225 0.615 ;
      RECT 2.61 0.255 4.225 0.425 ;
      RECT 2.61 0.425 2.78 0.84 ;
      RECT 1.615 0.84 2.78 1.01 ;
      RECT 1.615 1.01 1.785 2.735 ;
      RECT 1.615 0.575 1.865 0.84 ;
      RECT 1.005 2.905 2.125 3.075 ;
      RECT 1.955 1.855 2.125 2.905 ;
      RECT 1.955 1.685 3.23 1.855 ;
      RECT 2.975 1.855 3.23 2.355 ;
      RECT 3.005 1.455 3.23 1.685 ;
      RECT 3.005 1.125 3.545 1.455 ;
      RECT 1.005 1.82 1.445 2.905 ;
      RECT 1.275 1.13 1.445 1.82 ;
      RECT 1.055 0.35 1.445 1.13 ;
      RECT 8.765 1.78 8.995 2.12 ;
      RECT 8.765 1.45 9.16 1.78 ;
      RECT 12.635 1.27 13.695 1.6 ;
      RECT 12.545 1.82 12.875 2.86 ;
      RECT 12.635 1.6 12.875 1.82 ;
      RECT 12.635 0.35 12.885 1.27 ;
      RECT 0 -0.085 14.4 0.085 ;
      RECT 13.97 0.085 14.3 0.68 ;
      RECT 12.155 0.085 12.405 1.26 ;
      RECT 13.095 0.085 13.37 1.05 ;
      RECT 2.045 0.085 2.44 0.67 ;
      RECT 5.745 0.085 6.075 1.025 ;
      RECT 8.785 0.085 8.955 0.84 ;
      RECT 10.665 0.085 11.45 0.5 ;
      RECT 0.545 0.085 0.875 0.79 ;
      RECT 0 3.245 14.4 3.415 ;
      RECT 14.045 2.11 14.295 3.245 ;
      RECT 12.015 2.19 12.345 3.245 ;
      RECT 13.065 1.82 13.315 3.245 ;
      RECT 8.01 2.97 8.34 3.245 ;
      RECT 9.105 2.97 9.435 3.245 ;
      RECT 5.055 2.66 5.385 3.245 ;
      RECT 6.095 2.66 6.425 3.245 ;
      RECT 11.115 2.63 11.445 3.245 ;
      RECT 2.295 2.525 2.465 3.245 ;
      RECT 0.635 2.29 0.805 3.245 ;
  END
END scs8ls_dfbbn_2

MACRO scs8ls_dfbbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.24 1.47 8.57 1.74 ;
        RECT 7.28 1.74 8.57 1.8 ;
        RECT 7.28 1.8 8.515 1.91 ;
        RECT 7.28 1.91 7.45 2.905 ;
        RECT 6.04 2.905 7.45 3.075 ;
        RECT 6.04 2.335 6.21 2.905 ;
        RECT 5.16 2.165 6.21 2.335 ;
        RECT 5.16 2.335 5.33 2.905 ;
        RECT 4.36 2.905 5.33 3.075 ;
        RECT 4.36 1.655 4.53 2.905 ;
        RECT 4.23 1.41 4.56 1.655 ;
    END
    ANTENNAGATEAREA 0.47 ;
  END SETB

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.12 1.82 11.46 2.98 ;
        RECT 11.29 1.13 11.46 1.82 ;
        RECT 11.065 0.35 11.46 1.13 ;
    END
    ANTENNADIFFAREA 0.5189 ;
  END QN

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.235 0.98 10.58 1.65 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END RESETB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.96 1.825 2.29 2.155 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.18 0.805 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.525 0.35 12.86 2.98 ;
    END
    ANTENNADIFFAREA 0.519 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12.96 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12.96 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 9.755 1.21 9.925 1.38 ;
      RECT 5.435 1.21 5.605 1.38 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
    LAYER met1 ;
      RECT 5.375 1.365 5.665 1.41 ;
      RECT 5.375 1.225 9.985 1.365 ;
      RECT 9.695 1.365 9.985 1.41 ;
      RECT 5.375 1.18 5.665 1.225 ;
      RECT 9.695 1.18 9.985 1.225 ;
    LAYER li1 ;
      RECT 11.64 2.03 11.89 2.91 ;
      RECT 11.64 1.585 11.81 2.03 ;
      RECT 11.64 1.255 12.355 1.585 ;
      RECT 11.64 0.35 11.875 1.255 ;
      RECT 9.71 1.82 10.405 2.07 ;
      RECT 9.895 0.35 10.385 0.81 ;
      RECT 9.71 1.19 10.065 1.82 ;
      RECT 9.895 0.81 10.065 1.19 ;
      RECT 10.78 1.32 11.12 1.65 ;
      RECT 8.685 2.38 10.95 2.41 ;
      RECT 7.62 2.24 10.95 2.38 ;
      RECT 10.78 1.65 10.95 2.24 ;
      RECT 8.685 2.41 8.935 2.98 ;
      RECT 7.62 2.08 9.385 2.24 ;
      RECT 8.685 1.97 9.385 2.08 ;
      RECT 9.215 0.96 9.385 1.97 ;
      RECT 9.085 0.595 9.385 0.96 ;
      RECT 3.89 1.07 4.915 1.24 ;
      RECT 4.745 1.24 4.915 1.255 ;
      RECT 4.745 1.255 5.1 1.585 ;
      RECT 3.125 1.795 3.43 2.335 ;
      RECT 3.125 1.625 4.06 1.795 ;
      RECT 3.89 1.24 4.06 1.625 ;
      RECT 3.125 0.745 3.295 1.625 ;
      RECT 2.575 0.415 3.295 0.745 ;
      RECT 5.31 1.18 5.64 1.585 ;
      RECT 0.085 1.89 0.535 2.98 ;
      RECT 0.085 1.72 1.145 1.89 ;
      RECT 0.975 1.3 1.145 1.72 ;
      RECT 0.085 0.35 0.445 1.01 ;
      RECT 0.085 1.01 0.255 1.72 ;
      RECT 7.9 1.13 9.045 1.3 ;
      RECT 8.78 1.3 9.045 1.55 ;
      RECT 6.54 2.28 6.87 2.735 ;
      RECT 6.54 2.11 7.11 2.28 ;
      RECT 6.94 1.57 7.11 2.11 ;
      RECT 6.94 0.595 7.175 1.4 ;
      RECT 6.94 1.4 8.07 1.57 ;
      RECT 7.9 1.3 8.07 1.4 ;
      RECT 0 3.245 12.96 3.415 ;
      RECT 12.075 1.82 12.325 3.245 ;
      RECT 7.62 2.65 8.42 3.245 ;
      RECT 9.47 2.58 9.8 3.245 ;
      RECT 10.59 2.58 10.92 3.245 ;
      RECT 1.805 2.425 2.41 3.245 ;
      RECT 3.94 1.965 4.19 3.245 ;
      RECT 5.5 2.505 5.87 3.245 ;
      RECT 0.705 2.06 1.035 3.245 ;
      RECT 0 -0.085 12.96 0.085 ;
      RECT 12.055 0.085 12.305 0.81 ;
      RECT 10.565 0.085 10.895 0.81 ;
      RECT 6.19 0.67 6.43 1.085 ;
      RECT 6.06 0.085 6.43 0.67 ;
      RECT 0.615 0.085 0.945 1.01 ;
      RECT 1.655 0.085 1.905 1.065 ;
      RECT 3.56 0.085 4.155 0.56 ;
      RECT 8.085 0.085 8.415 0.96 ;
      RECT 4.415 0.425 4.825 0.56 ;
      RECT 4.415 0.255 5.84 0.425 ;
      RECT 5.51 0.425 5.84 0.67 ;
      RECT 2.58 2.295 2.955 2.755 ;
      RECT 2.785 1.085 2.955 2.295 ;
      RECT 2.085 0.915 2.955 1.085 ;
      RECT 2.085 0.605 2.335 0.915 ;
      RECT 1.315 1.255 2.615 1.585 ;
      RECT 1.315 1.585 1.565 2.98 ;
      RECT 1.315 1.13 1.485 1.255 ;
      RECT 1.125 0.35 1.485 1.13 ;
      RECT 8.585 0.425 8.915 0.96 ;
      RECT 8.585 0.255 9.725 0.425 ;
      RECT 9.555 0.425 9.725 1.02 ;
      RECT 5.85 1.255 6.18 1.585 ;
      RECT 3.465 0.9 3.72 1.455 ;
      RECT 4.7 1.995 4.95 2.735 ;
      RECT 4.7 1.825 6.02 1.995 ;
      RECT 5.85 1.585 6.02 1.825 ;
      RECT 5.85 1.01 6.02 1.255 ;
      RECT 5.085 0.9 6.02 1.01 ;
      RECT 3.465 0.84 6.02 0.9 ;
      RECT 3.465 0.73 5.335 0.84 ;
      RECT 5.015 0.595 5.335 0.73 ;
      RECT 6.6 0.255 7.67 0.425 ;
      RECT 7.345 0.425 7.67 1.23 ;
      RECT 6.44 1.61 6.77 1.94 ;
      RECT 6.6 0.425 6.77 1.61 ;
  END
END scs8ls_dfbbp_1

MACRO scs8ls_dfrbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 11.52 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.26 1.81 9.95 2.985 ;
        RECT 9.56 0.35 9.95 1.81 ;
    END
    ANTENNADIFFAREA 0.9515 LAYER met1 ;
    ANTENNADIFFAREA 0.9515 LAYER met2 ;
    ANTENNADIFFAREA 0.9515 LAYER met3 ;
    ANTENNADIFFAREA 0.9515 LAYER met4 ;
    ANTENNADIFFAREA 0.9515 LAYER met5 ;
  END QN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1 0.52 2.195 ;
    END
    ANTENNAGATEAREA 0.126 LAYER met1 ;
    ANTENNAGATEAREA 0.126 LAYER met2 ;
    ANTENNAGATEAREA 0.126 LAYER met3 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ;
    ANTENNAGATEAREA 0.126 LAYER met5 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.81 1.31 2.275 1.695 ;
        RECT 2.045 1.695 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.261 LAYER met1 ;
    ANTENNAGATEAREA 0.261 LAYER met2 ;
    ANTENNAGATEAREA 0.261 LAYER met3 ;
    ANTENNAGATEAREA 0.261 LAYER met4 ;
    ANTENNAGATEAREA 0.261 LAYER met5 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.065 0.35 11.435 1.13 ;
        RECT 11.265 1.13 11.435 1.82 ;
        RECT 11.075 1.82 11.435 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 LAYER met1 ;
    ANTENNADIFFAREA 0.5413 LAYER met2 ;
    ANTENNADIFFAREA 0.5413 LAYER met3 ;
    ANTENNADIFFAREA 0.5413 LAYER met4 ;
    ANTENNADIFFAREA 0.5413 LAYER met5 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.52 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.52 3.575 ;
    END
  END vpwr

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.055 1.965 8.065 2.105 ;
        RECT 1.055 2.105 1.345 2.15 ;
        RECT 1.055 1.92 1.345 1.965 ;
        RECT 5.375 2.105 5.665 2.15 ;
        RECT 7.775 2.105 8.065 2.15 ;
        RECT 5.375 1.92 5.665 1.965 ;
        RECT 7.775 1.92 8.065 1.965 ;
    END
    ANTENNAGATEAREA 0.378 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.956 LAYER met1 ;
    ANTENNAGATEAREA 0.378 LAYER met2 ;
    ANTENNAGATEAREA 0.378 LAYER met3 ;
    ANTENNAGATEAREA 0.378 LAYER met4 ;
    ANTENNAGATEAREA 0.378 LAYER met5 ;
  END RESETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 1.95 1.285 2.12 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 1.95 8.005 2.12 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 1.95 5.605 2.12 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
    LAYER li1 ;
      RECT 10.19 1.3 11.095 1.63 ;
      RECT 10.19 1.63 10.44 2.975 ;
      RECT 10.19 0.35 10.44 1.3 ;
      RECT 8.26 2.335 8.64 2.73 ;
      RECT 8.47 1.935 8.64 2.335 ;
      RECT 8.47 1.765 8.97 1.935 ;
      RECT 8.8 1.07 8.97 1.765 ;
      RECT 7.43 0.9 8.97 1.07 ;
      RECT 7.43 1.07 7.76 1.23 ;
      RECT 8.485 0.35 8.97 0.9 ;
      RECT 6.7 2.365 7.665 2.695 ;
      RECT 7.495 1.595 7.665 2.365 ;
      RECT 6.99 1.425 8.63 1.595 ;
      RECT 8.33 1.265 8.63 1.425 ;
      RECT 6.99 0.73 7.16 1.425 ;
      RECT 6.425 0.4 7.16 0.73 ;
      RECT 7.835 1.835 8.3 2.165 ;
      RECT 2.475 2.08 2.975 2.24 ;
      RECT 2.475 2.065 3 2.08 ;
      RECT 2.475 2.06 3.02 2.065 ;
      RECT 2.475 2.04 3.025 2.06 ;
      RECT 2.475 2.015 3.05 2.04 ;
      RECT 2.475 1.865 3.5 2.015 ;
      RECT 2.915 1.825 3.5 1.865 ;
      RECT 2.945 1.795 3.5 1.825 ;
      RECT 2.975 1.575 3.5 1.795 ;
      RECT 2.975 1.39 3.16 1.575 ;
      RECT 2.945 1.205 3.16 1.39 ;
      RECT 2.945 0.805 3.115 1.205 ;
      RECT 2.61 0.425 3.115 0.805 ;
      RECT 2.61 0.255 4.52 0.425 ;
      RECT 4.35 0.425 4.52 0.58 ;
      RECT 4.35 0.58 6.255 0.75 ;
      RECT 6.085 0.75 6.255 0.9 ;
      RECT 6.085 0.9 6.82 1.23 ;
      RECT 6.65 1.23 6.82 1.865 ;
      RECT 6.65 1.865 7.325 2.195 ;
      RECT 6.23 1.57 6.48 2.755 ;
      RECT 5.745 1.4 6.48 1.57 ;
      RECT 5.745 1.09 5.915 1.4 ;
      RECT 4.35 0.92 5.915 1.09 ;
      RECT 4.35 1.09 4.63 2.155 ;
      RECT 5.23 1.825 5.61 2.155 ;
      RECT 4.99 2.54 5.325 2.68 ;
      RECT 4.945 2.495 5.325 2.54 ;
      RECT 4.01 2.325 5.325 2.495 ;
      RECT 4.01 2.495 4.27 2.525 ;
      RECT 4.89 2.28 5.105 2.325 ;
      RECT 4.01 1.03 4.18 2.325 ;
      RECT 3.515 2.525 4.27 2.695 ;
      RECT 4.89 1.615 5.06 2.28 ;
      RECT 3.705 0.595 4.18 1.03 ;
      RECT 4.89 1.445 5.56 1.615 ;
      RECT 5.23 1.285 5.56 1.445 ;
      RECT 0.565 2.52 3.345 2.58 ;
      RECT 3.065 2.58 3.345 2.69 ;
      RECT 0.69 2.42 3.345 2.52 ;
      RECT 1.89 2.41 3.345 2.42 ;
      RECT 3.145 2.355 3.345 2.41 ;
      RECT 3.145 2.185 3.84 2.355 ;
      RECT 3.67 1.37 3.84 2.185 ;
      RECT 3.33 1.2 3.84 1.37 ;
      RECT 3.33 1.035 3.535 1.2 ;
      RECT 3.285 0.595 3.535 1.035 ;
      RECT 0.565 2.63 0.845 2.98 ;
      RECT 0.565 2.58 0.89 2.63 ;
      RECT 0.69 2.41 1.53 2.42 ;
      RECT 0.69 2.31 1.425 2.41 ;
      RECT 0.69 0.83 0.86 2.31 ;
      RECT 0.17 0.66 0.86 0.83 ;
      RECT 0.17 0.37 0.5 0.66 ;
      RECT 1.405 2.58 1.965 2.59 ;
      RECT 1.47 0.975 2.775 1.14 ;
      RECT 2.445 1.14 2.775 1.49 ;
      RECT 1.47 0.97 2.56 0.975 ;
      RECT 2.445 1.49 2.805 1.55 ;
      RECT 2.475 1.55 2.805 1.695 ;
      RECT 1.47 1.14 1.64 1.865 ;
      RECT 1.595 2.14 1.825 2.25 ;
      RECT 1.47 1.865 1.825 2.14 ;
      RECT 1.47 0.595 1.92 0.97 ;
      RECT 0 3.245 11.52 3.415 ;
      RECT 10.61 1.82 10.905 3.245 ;
      RECT 2.025 2.75 2.355 3.245 ;
      RECT 4.44 2.665 4.785 3.245 ;
      RECT 7.835 2.335 8.06 3.245 ;
      RECT 8.81 2.105 9.025 3.245 ;
      RECT 5.78 1.74 6.03 3.245 ;
      RECT 1.015 2.75 1.345 3.245 ;
      RECT 0.115 2.52 0.365 3.245 ;
      RECT 0 -0.085 11.52 0.085 ;
      RECT 10.645 0.085 10.895 1.13 ;
      RECT 1.03 0.085 1.28 0.83 ;
      RECT 2.09 0.085 2.42 0.8 ;
      RECT 4.995 0.085 5.325 0.41 ;
      RECT 7.535 0.085 7.995 0.68 ;
      RECT 9.14 0.085 9.39 1.13 ;
      RECT 1.03 1.13 1.3 2.14 ;
  END
END scs8ls_dfrbp_1

MACRO scs8ls_dfrbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 13.92 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.705 1.18 7.045 1.67 ;
    END
    ANTENNAGATEAREA 0.279 LAYER met1 ;
    ANTENNAGATEAREA 0.279 LAYER met2 ;
    ANTENNAGATEAREA 0.279 LAYER met3 ;
    ANTENNAGATEAREA 0.279 LAYER met4 ;
    ANTENNAGATEAREA 0.279 LAYER met5 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.81 0.515 1.57 ;
    END
    ANTENNAGATEAREA 0.126 LAYER met1 ;
    ANTENNAGATEAREA 0.126 LAYER met2 ;
    ANTENNAGATEAREA 0.126 LAYER met3 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ;
    ANTENNAGATEAREA 0.126 LAYER met5 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.195 0.77 11.875 1.32 ;
        RECT 10.895 1.32 11.875 1.41 ;
        RECT 11.195 0.35 11.455 0.77 ;
        RECT 10.895 1.41 11.725 1.54 ;
        RECT 10.895 1.54 11.065 2.9 ;
    END
    ANTENNADIFFAREA 0.5432 LAYER met1 ;
    ANTENNADIFFAREA 0.5432 LAYER met2 ;
    ANTENNADIFFAREA 0.5432 LAYER met3 ;
    ANTENNADIFFAREA 0.5432 LAYER met4 ;
    ANTENNADIFFAREA 0.5432 LAYER met5 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.06 0.33 13.39 1.13 ;
        RECT 13.135 1.13 13.305 1.82 ;
        RECT 12.975 1.82 13.305 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 LAYER met1 ;
    ANTENNADIFFAREA 0.5432 LAYER met2 ;
    ANTENNADIFFAREA 0.5432 LAYER met3 ;
    ANTENNADIFFAREA 0.5432 LAYER met4 ;
    ANTENNADIFFAREA 0.5432 LAYER met5 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.92 3.575 ;
    END
  END vpwr

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.055 1.595 9.985 1.735 ;
        RECT 2.495 1.735 2.785 1.78 ;
        RECT 2.495 1.55 2.785 1.595 ;
        RECT 1.055 1.735 1.345 1.78 ;
        RECT 9.695 1.735 9.985 1.78 ;
        RECT 1.055 1.55 1.345 1.595 ;
        RECT 9.695 1.55 9.985 1.595 ;
    END
    ANTENNAGATEAREA 0.378 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3 LAYER met1 ;
    ANTENNAGATEAREA 0.378 LAYER met2 ;
    ANTENNAGATEAREA 0.378 LAYER met3 ;
    ANTENNAGATEAREA 0.378 LAYER met4 ;
    ANTENNAGATEAREA 0.378 LAYER met5 ;
  END RESETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 1.58 9.925 1.75 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 1.58 2.725 1.75 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 1.58 1.285 1.75 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
    LAYER li1 ;
      RECT 0 3.245 13.92 3.415 ;
      RECT 13.475 1.82 13.805 3.245 ;
      RECT 12.475 1.82 12.805 3.245 ;
      RECT 11.265 1.74 11.595 3.245 ;
      RECT 0.115 2.965 1.435 3.245 ;
      RECT 5.99 2.765 6.5 3.245 ;
      RECT 2.945 2.625 3.195 3.245 ;
      RECT 9.265 2.29 9.625 3.245 ;
      RECT 10.365 2.29 10.695 3.245 ;
      RECT 0.115 1.94 0.51 2.965 ;
      RECT 0 -0.085 13.92 0.085 ;
      RECT 13.56 0.085 13.82 1.13 ;
      RECT 11.625 0.085 11.965 0.6 ;
      RECT 12.63 0.085 12.88 1.13 ;
      RECT 1.145 0.085 1.475 0.81 ;
      RECT 2.205 0.085 2.535 0.78 ;
      RECT 5.605 0.085 5.855 0.49 ;
      RECT 9.415 0.085 9.745 0.72 ;
      RECT 10.845 0.085 11.015 1.1 ;
      RECT 6.705 2.17 7.035 2.255 ;
      RECT 6.095 1.84 7.505 2.17 ;
      RECT 6.365 0.635 6.96 0.965 ;
      RECT 6.095 1.67 6.265 1.84 ;
      RECT 5.595 1.34 6.535 1.67 ;
      RECT 6.365 0.965 6.535 1.34 ;
      RECT 9.83 2.12 10.16 2.385 ;
      RECT 9.065 1.95 10.675 2.12 ;
      RECT 9.065 1.455 9.33 1.95 ;
      RECT 10.505 0.765 10.675 1.95 ;
      RECT 10.205 0.35 10.675 0.765 ;
      RECT 1.605 2.905 2.775 3.075 ;
      RECT 1.605 2.795 1.775 2.905 ;
      RECT 2.605 2.455 2.775 2.905 ;
      RECT 0.68 2.625 1.775 2.795 ;
      RECT 2.605 2.285 3.535 2.455 ;
      RECT 0.68 1.95 1.01 2.625 ;
      RECT 3.365 2.455 3.535 2.905 ;
      RECT 0.685 0.64 0.855 1.95 ;
      RECT 3.365 2.905 4.46 3.075 ;
      RECT 0.325 0.39 0.855 0.64 ;
      RECT 4.29 2.815 4.46 2.905 ;
      RECT 4.29 2.485 4.96 2.815 ;
      RECT 4.29 2.41 4.475 2.485 ;
      RECT 4.305 1.105 4.475 2.41 ;
      RECT 3.345 0.935 4.475 1.105 ;
      RECT 3.345 1.105 3.715 1.385 ;
      RECT 9.54 1.45 9.955 1.78 ;
      RECT 7.555 0.765 7.725 1.185 ;
      RECT 7.555 0.595 9.235 0.765 ;
      RECT 8.985 0.35 9.235 0.595 ;
      RECT 11.895 1.74 12.305 2.78 ;
      RECT 12.135 1.63 12.305 1.74 ;
      RECT 12.135 1.3 12.965 1.63 ;
      RECT 12.135 0.35 12.43 1.3 ;
      RECT 4.645 0.765 4.895 1.6 ;
      RECT 3.045 0.595 4.895 0.765 ;
      RECT 2.185 2.115 2.435 2.735 ;
      RECT 1.825 1.945 4.12 2.115 ;
      RECT 3.79 2.115 4.12 2.735 ;
      RECT 3.885 1.61 4.12 1.945 ;
      RECT 1.825 1.47 2.155 1.945 ;
      RECT 3.885 1.275 4.135 1.61 ;
      RECT 2.385 1.445 2.755 1.775 ;
      RECT 1.025 1.45 1.315 1.78 ;
      RECT 5.425 2.425 7.505 2.595 ;
      RECT 7.315 2.595 7.505 2.905 ;
      RECT 7.315 2.905 8.22 3.075 ;
      RECT 8.05 1.605 8.22 2.905 ;
      RECT 8.05 1.275 8.555 1.605 ;
      RECT 5.425 2.595 5.785 2.98 ;
      RECT 5.425 2.24 5.785 2.425 ;
      RECT 4.645 1.91 5.785 2.24 ;
      RECT 5.095 1.84 5.785 1.91 ;
      RECT 5.095 1 5.425 1.84 ;
      RECT 8.39 2.095 8.64 2.385 ;
      RECT 8.39 1.925 8.895 2.095 ;
      RECT 8.725 1.265 8.895 1.925 ;
      RECT 8.725 1.105 10.335 1.265 ;
      RECT 7.905 0.935 10.335 1.105 ;
      RECT 6.025 0.255 8.78 0.425 ;
      RECT 7.215 0.425 7.385 1.355 ;
      RECT 7.215 1.355 7.88 1.525 ;
      RECT 7.71 1.525 7.88 2.735 ;
      RECT 1.485 2.285 1.97 2.455 ;
      RECT 1.485 1.185 1.655 2.285 ;
      RECT 1.485 1.015 3.095 1.185 ;
      RECT 2.925 1.185 3.095 1.555 ;
      RECT 1.645 0.465 1.975 1.015 ;
      RECT 2.705 0.425 2.875 1.015 ;
      RECT 2.925 1.555 3.255 1.775 ;
      RECT 2.705 0.255 5.235 0.425 ;
      RECT 5.065 0.425 5.235 0.66 ;
      RECT 5.065 0.66 6.195 0.83 ;
      RECT 6.025 0.425 6.195 0.66 ;
  END
END scs8ls_dfrbp_2

MACRO scs8ls_dfrtn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 11.04 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.96 0.37 2.15 ;
    END
    ANTENNAGATEAREA 0.126 LAYER met1 ;
    ANTENNAGATEAREA 0.126 LAYER met2 ;
    ANTENNAGATEAREA 0.126 LAYER met3 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ;
    ANTENNAGATEAREA 0.126 LAYER met5 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.605 1.82 10.955 2.98 ;
        RECT 10.785 1.15 10.955 1.82 ;
        RECT 10.59 0.44 10.955 1.15 ;
    END
    ANTENNADIFFAREA 0.5338 LAYER met1 ;
    ANTENNADIFFAREA 0.5338 LAYER met2 ;
    ANTENNADIFFAREA 0.5338 LAYER met3 ;
    ANTENNADIFFAREA 0.5338 LAYER met4 ;
    ANTENNADIFFAREA 0.5338 LAYER met5 ;
  END Q

  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.455 1.18 1.765 1.65 ;
    END
    ANTENNAGATEAREA 0.261 LAYER met1 ;
    ANTENNAGATEAREA 0.261 LAYER met2 ;
    ANTENNAGATEAREA 0.261 LAYER met3 ;
    ANTENNAGATEAREA 0.261 LAYER met4 ;
    ANTENNAGATEAREA 0.261 LAYER met5 ;
  END CLKN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.04 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.04 3.575 ;
    END
  END vpwr

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.055 1.595 8.545 1.735 ;
        RECT 1.055 1.735 1.345 1.78 ;
        RECT 4.895 1.735 5.185 1.78 ;
        RECT 8.255 1.735 8.545 1.78 ;
        RECT 1.055 1.55 1.345 1.595 ;
        RECT 4.895 1.55 5.185 1.595 ;
        RECT 8.255 1.55 8.545 1.595 ;
    END
    ANTENNAGATEAREA 0.378 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 5.292 LAYER met1 ;
    ANTENNAGATEAREA 0.378 LAYER met2 ;
    ANTENNAGATEAREA 0.378 LAYER met3 ;
    ANTENNAGATEAREA 0.378 LAYER met4 ;
    ANTENNAGATEAREA 0.378 LAYER met5 ;
  END RESETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 1.58 8.485 1.75 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 1.58 5.125 1.75 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 1.58 1.285 1.75 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
    LAYER li1 ;
      RECT 0.54 2.18 3.42 2.35 ;
      RECT 3.17 2.35 3.42 2.735 ;
      RECT 2.335 0.725 2.505 2.18 ;
      RECT 2.335 0.705 2.535 0.725 ;
      RECT 2.335 0.685 2.55 0.705 ;
      RECT 2.335 0.655 2.575 0.685 ;
      RECT 2.335 0.625 3.365 0.655 ;
      RECT 3.115 0.655 3.365 1.075 ;
      RECT 2.355 0.605 3.365 0.625 ;
      RECT 2.37 0.595 3.365 0.605 ;
      RECT 2.395 0.565 3.365 0.595 ;
      RECT 2.41 0.545 3.365 0.565 ;
      RECT 2.415 0.525 3.365 0.545 ;
      RECT 2.44 0.485 3.365 0.525 ;
      RECT 0.64 2.35 0.87 2.98 ;
      RECT 0.54 0.79 0.71 2.18 ;
      RECT 0.145 0.35 0.71 0.79 ;
      RECT 0 -0.085 11.04 0.085 ;
      RECT 1.045 0.085 1.295 0.81 ;
      RECT 2.02 0.085 2.255 0.465 ;
      RECT 5.025 0.085 5.355 0.62 ;
      RECT 8.115 0.085 8.555 0.905 ;
      RECT 10.16 0.085 10.41 1.13 ;
      RECT 8.285 1.465 8.71 1.795 ;
      RECT 3.62 2.18 4.075 2.735 ;
      RECT 3.875 2.14 4.075 2.18 ;
      RECT 3.875 1.97 5.695 2.14 ;
      RECT 4.97 2.14 5.3 2.735 ;
      RECT 5.335 1.47 5.695 1.97 ;
      RECT 3.875 0.635 4.075 1.97 ;
      RECT 8.68 2.335 9.01 2.98 ;
      RECT 8.07 2.135 9.05 2.335 ;
      RECT 8.07 1.965 9.56 2.135 ;
      RECT 9.39 0.955 9.56 1.965 ;
      RECT 9.045 0.575 9.56 0.955 ;
      RECT 6.87 2.705 7.6 2.865 ;
      RECT 6.87 2.535 7.9 2.705 ;
      RECT 7.73 1.295 7.9 2.535 ;
      RECT 7.73 1.125 9.22 1.295 ;
      RECT 8.92 1.295 9.22 1.795 ;
      RECT 7.73 0.955 7.9 1.125 ;
      RECT 6.705 0.625 7.9 0.955 ;
      RECT 1.515 1.82 2.165 2.01 ;
      RECT 1.935 1.01 2.165 1.82 ;
      RECT 1.475 0.665 2.165 1.01 ;
      RECT 1.475 0.35 1.805 0.665 ;
      RECT 0 3.245 11.04 3.415 ;
      RECT 0.11 2.52 0.44 3.245 ;
      RECT 1.04 2.52 1.37 3.245 ;
      RECT 2.07 2.52 2.4 3.245 ;
      RECT 8.14 2.52 8.47 3.245 ;
      RECT 9.21 2.52 9.46 3.245 ;
      RECT 5.49 2.36 5.82 3.245 ;
      RECT 4.46 2.31 4.79 3.245 ;
      RECT 10.15 2.1 10.4 3.245 ;
      RECT 7.31 1.8 7.56 2.365 ;
      RECT 6.205 1.63 7.56 1.8 ;
      RECT 6.205 1.47 6.51 1.63 ;
      RECT 0.88 1.245 1.285 1.78 ;
      RECT 4.855 1.47 5.155 1.8 ;
      RECT 5.99 2.14 6.7 2.98 ;
      RECT 5.865 1.97 6.7 2.14 ;
      RECT 5.865 1.3 6.035 1.97 ;
      RECT 4.275 1.13 6.195 1.3 ;
      RECT 4.275 1.3 4.655 1.775 ;
      RECT 5.865 0.595 6.195 1.13 ;
      RECT 6.75 1.295 7.42 1.455 ;
      RECT 6.365 1.125 7.42 1.295 ;
      RECT 6.365 0.425 6.535 1.125 ;
      RECT 5.525 0.255 6.535 0.425 ;
      RECT 5.525 0.425 5.695 0.79 ;
      RECT 4.685 0.79 5.695 0.96 ;
      RECT 4.685 0.465 4.855 0.79 ;
      RECT 3.535 0.255 4.855 0.465 ;
      RECT 3.535 0.465 3.705 1.245 ;
      RECT 2.675 1.245 3.705 2.01 ;
      RECT 2.675 0.825 2.94 1.245 ;
      RECT 9.73 1.32 10.615 1.65 ;
      RECT 9.65 2.305 9.98 2.98 ;
      RECT 9.73 1.65 9.98 2.305 ;
      RECT 9.73 0.53 9.98 1.32 ;
  END
END scs8ls_dfrtn_1

MACRO scs8ls_dfrtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 11.04 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1 0.515 2.17 ;
    END
    ANTENNAGATEAREA 0.126 LAYER met1 ;
    ANTENNAGATEAREA 0.126 LAYER met2 ;
    ANTENNAGATEAREA 0.126 LAYER met3 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ;
    ANTENNAGATEAREA 0.126 LAYER met5 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.795 1.31 2.275 1.775 ;
        RECT 2.045 1.775 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.261 LAYER met1 ;
    ANTENNAGATEAREA 0.261 LAYER met2 ;
    ANTENNAGATEAREA 0.261 LAYER met3 ;
    ANTENNAGATEAREA 0.261 LAYER met4 ;
    ANTENNAGATEAREA 0.261 LAYER met5 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.725 1.885 10.425 2.98 ;
        RECT 10.165 1.13 10.425 1.885 ;
        RECT 10.165 0.35 10.495 1.13 ;
    END
    ANTENNADIFFAREA 0.5917 LAYER met1 ;
    ANTENNADIFFAREA 0.5917 LAYER met2 ;
    ANTENNADIFFAREA 0.5917 LAYER met3 ;
    ANTENNADIFFAREA 0.5917 LAYER met4 ;
    ANTENNADIFFAREA 0.5917 LAYER met5 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.04 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.04 3.575 ;
    END
  END vpwr

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.055 1.965 8.065 2.105 ;
        RECT 1.055 2.105 1.345 2.15 ;
        RECT 1.055 1.92 1.345 1.965 ;
        RECT 4.895 2.105 5.185 2.15 ;
        RECT 7.775 2.105 8.065 2.15 ;
        RECT 4.895 1.92 5.185 1.965 ;
        RECT 7.775 1.92 8.065 1.965 ;
    END
    ANTENNAGATEAREA 0.378 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.956 LAYER met1 ;
    ANTENNAGATEAREA 0.378 LAYER met2 ;
    ANTENNAGATEAREA 0.378 LAYER met3 ;
    ANTENNAGATEAREA 0.378 LAYER met4 ;
    ANTENNAGATEAREA 0.378 LAYER met5 ;
  END RESETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.835 1.95 8.005 2.12 ;
      RECT 4.955 1.95 5.125 2.12 ;
      RECT 1.115 1.95 1.285 2.12 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
    LAYER li1 ;
      RECT 10.675 0.085 10.925 1.13 ;
      RECT 0 -0.085 11.04 0.085 ;
      RECT 4.915 0.085 5.31 0.395 ;
      RECT 7.745 0.085 8.075 0.845 ;
      RECT 9.175 0.085 9.425 0.845 ;
      RECT 1.03 0.085 1.28 0.83 ;
      RECT 2.06 0.085 2.39 0.8 ;
      RECT 4.615 2.32 5.25 2.4 ;
      RECT 4.615 1.575 4.785 2.32 ;
      RECT 3.46 2.57 4.215 2.725 ;
      RECT 3.93 1.05 4.1 2.4 ;
      RECT 4.615 1.245 5.65 1.575 ;
      RECT 3.625 0.67 4.1 1.05 ;
      RECT 3.46 2.495 5.25 2.57 ;
      RECT 3.93 2.4 5.25 2.495 ;
      RECT 10.595 1.82 10.925 3.245 ;
      RECT 0 3.245 11.04 3.415 ;
      RECT 1.985 2.74 2.315 3.245 ;
      RECT 7.805 2.445 8.135 3.245 ;
      RECT 8.855 2.195 9.185 3.245 ;
      RECT 5.48 1.745 5.81 3.245 ;
      RECT 4.385 2.74 4.715 3.245 ;
      RECT 0.105 2.52 0.355 3.245 ;
      RECT 0.98 2.73 1.31 3.245 ;
      RECT 6.965 1.345 7.295 2.305 ;
      RECT 6.69 1.015 7.42 1.345 ;
      RECT 7.25 0.425 7.42 1.015 ;
      RECT 5.48 0.255 7.42 0.425 ;
      RECT 5.48 0.425 5.65 0.565 ;
      RECT 4.27 0.5 4.44 0.565 ;
      RECT 2.56 0.33 4.44 0.5 ;
      RECT 2.56 0.5 3.035 0.805 ;
      RECT 2.865 0.805 3.035 1.195 ;
      RECT 2.865 1.195 3.115 1.345 ;
      RECT 2.945 1.345 3.115 1.56 ;
      RECT 2.945 1.56 3.42 1.82 ;
      RECT 2.9 1.82 3.42 1.865 ;
      RECT 2.445 1.865 3.42 1.985 ;
      RECT 2.445 1.985 3.06 2.035 ;
      RECT 2.445 2.035 2.775 2.205 ;
      RECT 4.27 0.565 5.65 0.735 ;
      RECT 1.405 2.56 3.29 2.57 ;
      RECT 3.01 2.57 3.29 2.725 ;
      RECT 1.835 2.405 3.29 2.41 ;
      RECT 1.85 2.4 3.29 2.405 ;
      RECT 1.87 2.39 3.29 2.4 ;
      RECT 1.895 2.375 3.29 2.39 ;
      RECT 3.01 2.37 3.29 2.375 ;
      RECT 3.01 2.325 3.335 2.37 ;
      RECT 3.01 2.205 3.76 2.325 ;
      RECT 3.185 2.155 3.76 2.205 ;
      RECT 3.59 1.39 3.76 2.155 ;
      RECT 3.285 1.22 3.76 1.39 ;
      RECT 3.285 1.045 3.455 1.22 ;
      RECT 3.205 0.67 3.455 1.045 ;
      RECT 0.555 2.52 3.29 2.56 ;
      RECT 0.685 2.41 3.29 2.52 ;
      RECT 0.555 2.56 0.86 2.605 ;
      RECT 0.685 0.83 0.855 2.31 ;
      RECT 0.555 2.605 0.835 2.64 ;
      RECT 0.13 0.66 0.855 0.83 ;
      RECT 0.555 2.64 0.81 2.98 ;
      RECT 0.13 0.37 0.46 0.66 ;
      RECT 0.685 2.39 1.53 2.41 ;
      RECT 0.685 2.375 1.51 2.39 ;
      RECT 0.685 2.36 1.49 2.375 ;
      RECT 0.685 2.335 1.465 2.36 ;
      RECT 0.685 2.31 1.435 2.335 ;
      RECT 1.435 2.59 1.86 2.61 ;
      RECT 1.435 2.585 1.89 2.59 ;
      RECT 1.405 2.58 1.89 2.585 ;
      RECT 1.405 2.575 1.91 2.58 ;
      RECT 1.405 2.57 1.925 2.575 ;
      RECT 9.385 1.385 9.935 1.715 ;
      RECT 9.605 0.35 9.935 1.385 ;
      RECT 9.385 1.715 9.555 2.905 ;
      RECT 1.025 1.13 1.285 2.14 ;
      RECT 1.455 0.975 2.695 1.14 ;
      RECT 2.445 1.14 2.695 1.49 ;
      RECT 1.455 0.97 2.505 0.975 ;
      RECT 2.445 1.49 2.775 1.695 ;
      RECT 1.615 2.205 1.785 2.24 ;
      RECT 1.455 1.14 1.625 1.945 ;
      RECT 1.615 2.14 1.865 2.205 ;
      RECT 1.455 1.945 1.865 2.14 ;
      RECT 1.455 0.35 1.84 0.97 ;
      RECT 4.27 1.075 4.445 2.125 ;
      RECT 5.82 1.075 6.15 1.13 ;
      RECT 5.82 0.665 6.15 0.905 ;
      RECT 5.98 1.13 6.15 1.865 ;
      RECT 5.98 1.865 6.31 2.755 ;
      RECT 4.27 0.905 6.15 1.075 ;
      RECT 4.955 1.795 5.285 2.15 ;
      RECT 8.32 2.445 8.685 2.905 ;
      RECT 8.515 2.025 8.685 2.445 ;
      RECT 8.515 1.855 9.19 2.025 ;
      RECT 9.02 1.185 9.19 1.855 ;
      RECT 7.59 1.015 9.19 1.185 ;
      RECT 7.59 1.185 7.92 1.345 ;
      RECT 8.615 0.385 8.945 1.015 ;
      RECT 6.48 2.475 7.635 2.805 ;
      RECT 6.48 1.685 6.65 2.475 ;
      RECT 7.465 1.685 7.635 2.475 ;
      RECT 6.32 1.515 6.65 1.685 ;
      RECT 7.465 1.515 8.85 1.685 ;
      RECT 6.32 0.845 6.49 1.515 ;
      RECT 8.52 1.355 8.85 1.515 ;
      RECT 6.32 0.595 7.08 0.845 ;
      RECT 7.805 1.92 8.345 2.255 ;
  END
END scs8ls_dfrtp_1

MACRO scs8ls_dfrtp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 11.52 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.65 0.35 10.98 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 LAYER met1 ;
    ANTENNADIFFAREA 0.5432 LAYER met2 ;
    ANTENNADIFFAREA 0.5432 LAYER met3 ;
    ANTENNADIFFAREA 0.5432 LAYER met4 ;
    ANTENNADIFFAREA 0.5432 LAYER met5 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.795 1.32 2.275 1.73 ;
        RECT 2.045 1.73 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.261 LAYER met1 ;
    ANTENNAGATEAREA 0.261 LAYER met2 ;
    ANTENNAGATEAREA 0.261 LAYER met3 ;
    ANTENNAGATEAREA 0.261 LAYER met4 ;
    ANTENNAGATEAREA 0.261 LAYER met5 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1 0.495 2.17 ;
    END
    ANTENNAGATEAREA 0.126 LAYER met1 ;
    ANTENNAGATEAREA 0.126 LAYER met2 ;
    ANTENNAGATEAREA 0.126 LAYER met3 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ;
    ANTENNAGATEAREA 0.126 LAYER met5 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.52 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.52 3.575 ;
    END
  END vpwr

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.055 1.965 8.065 2.105 ;
        RECT 1.055 2.105 1.345 2.15 ;
        RECT 1.055 1.92 1.345 1.965 ;
        RECT 4.895 2.105 5.185 2.15 ;
        RECT 7.775 2.105 8.065 2.15 ;
        RECT 4.895 1.92 5.185 1.965 ;
        RECT 7.775 1.92 8.065 1.965 ;
    END
    ANTENNAGATEAREA 0.378 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.956 LAYER met1 ;
    ANTENNAGATEAREA 0.378 LAYER met2 ;
    ANTENNAGATEAREA 0.378 LAYER met3 ;
    ANTENNAGATEAREA 0.378 LAYER met4 ;
    ANTENNAGATEAREA 0.378 LAYER met5 ;
  END RESETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 1.95 8.005 2.12 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 1.95 5.125 2.12 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 1.95 1.285 2.12 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
    LAYER li1 ;
      RECT 1.005 1.14 1.285 2.15 ;
      RECT 7.805 1.92 8.395 2.275 ;
      RECT 2.53 2.23 2.775 2.275 ;
      RECT 2.515 2.205 2.775 2.23 ;
      RECT 2.515 2.08 2.94 2.205 ;
      RECT 2.515 2.035 3.01 2.08 ;
      RECT 2.515 1.985 3.095 2.035 ;
      RECT 2.515 1.945 3.425 1.985 ;
      RECT 2.81 1.9 3.425 1.945 ;
      RECT 2.865 1.625 3.425 1.9 ;
      RECT 2.865 0.805 3.07 1.625 ;
      RECT 2.595 0.5 3.07 0.805 ;
      RECT 2.595 0.33 4.475 0.5 ;
      RECT 4.305 0.5 4.475 0.615 ;
      RECT 4.305 0.615 5.685 0.785 ;
      RECT 5.515 0.425 5.685 0.615 ;
      RECT 5.515 0.255 7.455 0.425 ;
      RECT 7.285 0.425 7.455 1.015 ;
      RECT 6.725 1.015 7.455 1.345 ;
      RECT 6.955 1.345 7.285 2.305 ;
      RECT 6.015 1.855 6.345 2.755 ;
      RECT 6.015 1.13 6.185 1.855 ;
      RECT 5.855 1.125 6.185 1.13 ;
      RECT 4.275 0.955 6.185 1.125 ;
      RECT 4.275 1.125 4.445 2.125 ;
      RECT 5.855 0.595 6.185 0.955 ;
      RECT 0 3.245 11.52 3.415 ;
      RECT 11.155 1.82 11.405 3.245 ;
      RECT 1.955 2.74 2.285 3.245 ;
      RECT 4.42 2.74 4.75 3.245 ;
      RECT 7.795 2.445 8.125 3.245 ;
      RECT 9.09 2.445 9.42 3.245 ;
      RECT 10.15 1.82 10.48 3.245 ;
      RECT 5.515 1.745 5.845 3.245 ;
      RECT 1.015 2.73 1.345 3.245 ;
      RECT 0.105 2.52 0.435 3.245 ;
      RECT 3.495 2.57 4.25 2.75 ;
      RECT 3.495 2.525 5.285 2.57 ;
      RECT 3.935 2.4 5.285 2.525 ;
      RECT 4.615 2.32 5.285 2.4 ;
      RECT 3.935 1.05 4.105 2.4 ;
      RECT 4.615 1.575 4.785 2.32 ;
      RECT 3.66 0.67 4.105 1.05 ;
      RECT 4.615 1.295 5.685 1.575 ;
      RECT 9.59 2.03 9.92 2.905 ;
      RECT 9.66 1.63 9.92 2.03 ;
      RECT 9.66 1.3 10.19 1.63 ;
      RECT 9.66 0.35 9.99 1.3 ;
      RECT 4.955 1.795 5.285 2.15 ;
      RECT 0.635 2.52 3.325 2.56 ;
      RECT 1.405 2.56 3.325 2.57 ;
      RECT 0.665 2.445 3.325 2.52 ;
      RECT 2.33 2.57 3.325 2.575 ;
      RECT 0.665 2.44 2.485 2.445 ;
      RECT 2.945 2.4 3.325 2.445 ;
      RECT 2.345 2.575 3.325 2.58 ;
      RECT 0.665 2.435 2.47 2.44 ;
      RECT 2.945 2.375 3.37 2.4 ;
      RECT 2.355 2.58 3.325 2.585 ;
      RECT 0.665 2.43 2.46 2.435 ;
      RECT 3.11 2.355 3.37 2.375 ;
      RECT 2.365 2.585 3.325 2.59 ;
      RECT 0.665 2.42 2.44 2.43 ;
      RECT 3.11 2.23 3.765 2.355 ;
      RECT 2.375 2.59 3.325 2.595 ;
      RECT 0.665 2.405 2.42 2.42 ;
      RECT 3.2 2.185 3.765 2.23 ;
      RECT 2.39 2.595 3.325 2.605 ;
      RECT 0.665 2.395 2.405 2.405 ;
      RECT 3.595 1.39 3.765 2.185 ;
      RECT 2.405 2.605 3.325 2.615 ;
      RECT 0.665 2.38 2.385 2.395 ;
      RECT 3.32 1.22 3.765 1.39 ;
      RECT 3.045 2.615 3.325 2.725 ;
      RECT 0.665 2.355 2.36 2.38 ;
      RECT 3.32 1.045 3.49 1.22 ;
      RECT 0.665 2.33 2.34 2.355 ;
      RECT 3.24 0.67 3.49 1.045 ;
      RECT 0.635 2.63 0.835 2.98 ;
      RECT 0.635 2.605 0.87 2.63 ;
      RECT 0.635 2.56 0.89 2.605 ;
      RECT 0.665 0.83 0.835 2.33 ;
      RECT 0.13 0.66 0.835 0.83 ;
      RECT 0.13 0.37 0.46 0.66 ;
      RECT 6.515 2.475 7.625 2.805 ;
      RECT 7.455 1.73 7.625 2.475 ;
      RECT 6.515 1.685 6.685 2.475 ;
      RECT 7.455 1.56 9.035 1.73 ;
      RECT 6.355 1.515 6.685 1.685 ;
      RECT 8.705 1.73 9.035 1.89 ;
      RECT 6.355 0.845 6.525 1.515 ;
      RECT 6.355 0.595 7.115 0.845 ;
      RECT 8.295 2.445 8.885 2.775 ;
      RECT 8.715 2.275 8.885 2.445 ;
      RECT 8.715 2.105 9.375 2.275 ;
      RECT 9.205 1.39 9.375 2.105 ;
      RECT 7.625 1.22 9.375 1.39 ;
      RECT 7.625 1.06 7.955 1.22 ;
      RECT 8.68 0.385 9.01 1.22 ;
      RECT 0 -0.085 11.52 0.085 ;
      RECT 11.16 0.085 11.41 1.13 ;
      RECT 1.005 0.085 1.285 0.83 ;
      RECT 2.095 0.085 2.425 0.8 ;
      RECT 4.92 0.085 5.345 0.445 ;
      RECT 7.77 0.085 8.19 0.715 ;
      RECT 9.23 0.085 9.48 1.05 ;
      RECT 10.22 0.085 10.47 1.13 ;
      RECT 1.455 0.975 2.685 1.15 ;
      RECT 2.445 1.15 2.685 1.55 ;
      RECT 1.455 0.97 2.54 0.975 ;
      RECT 2.515 1.55 2.685 1.775 ;
      RECT 1.455 1.15 1.625 1.9 ;
      RECT 1.455 1.9 1.865 2.16 ;
      RECT 1.455 0.35 1.875 0.97 ;
  END
END scs8ls_dfrtp_2

MACRO scs8ls_dfrtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.41 1.61 13.315 1.78 ;
        RECT 12.41 1.78 12.74 1.8 ;
        RECT 12.575 1.27 13.315 1.61 ;
        RECT 11.035 1.8 12.74 1.97 ;
        RECT 12.575 1.13 12.825 1.27 ;
        RECT 11.035 1.97 11.365 2.98 ;
        RECT 12.41 1.97 12.74 2.98 ;
        RECT 11.595 0.88 12.825 1.13 ;
        RECT 11.595 0.365 11.91 0.88 ;
        RECT 12.575 0.35 12.825 0.88 ;
    END
    ANTENNADIFFAREA 1.2071 LAYER met1 ;
    ANTENNADIFFAREA 1.2071 LAYER met2 ;
    ANTENNADIFFAREA 1.2071 LAYER met3 ;
    ANTENNADIFFAREA 1.2071 LAYER met4 ;
    ANTENNADIFFAREA 1.2071 LAYER met5 ;
  END Q

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.845 1.64 2.275 1.775 ;
        RECT 2.045 1.775 2.275 1.78 ;
        RECT 1.795 1.31 2.275 1.64 ;
    END
    ANTENNAGATEAREA 0.261 LAYER met1 ;
    ANTENNAGATEAREA 0.261 LAYER met2 ;
    ANTENNAGATEAREA 0.261 LAYER met3 ;
    ANTENNAGATEAREA 0.261 LAYER met4 ;
    ANTENNAGATEAREA 0.261 LAYER met5 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1 0.515 2.18 ;
    END
    ANTENNAGATEAREA 0.126 LAYER met1 ;
    ANTENNAGATEAREA 0.126 LAYER met2 ;
    ANTENNAGATEAREA 0.126 LAYER met3 ;
    ANTENNAGATEAREA 0.126 LAYER met4 ;
    ANTENNAGATEAREA 0.126 LAYER met5 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.44 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.44 3.575 ;
    END
  END vpwr

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.055 1.965 9.025 2.105 ;
        RECT 1.055 2.105 1.345 2.15 ;
        RECT 1.055 1.92 1.345 1.965 ;
        RECT 5.375 2.105 5.665 2.15 ;
        RECT 8.735 2.105 9.025 2.15 ;
        RECT 5.375 1.92 5.665 1.965 ;
        RECT 8.735 1.92 9.025 1.965 ;
    END
    ANTENNAGATEAREA 0.378 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 5.628 LAYER met1 ;
    ANTENNAGATEAREA 0.378 LAYER met2 ;
    ANTENNAGATEAREA 0.378 LAYER met3 ;
    ANTENNAGATEAREA 0.378 LAYER met4 ;
    ANTENNAGATEAREA 0.378 LAYER met5 ;
  END RESETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 1.95 8.965 2.12 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 1.95 5.605 2.12 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 1.95 1.285 2.12 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
    LAYER li1 ;
      RECT 5.395 2.405 6.955 2.575 ;
      RECT 5.395 2.29 5.725 2.405 ;
      RECT 6.785 1.59 6.955 2.405 ;
      RECT 6.495 1.26 6.955 1.59 ;
      RECT 3.48 2.57 4.23 2.755 ;
      RECT 3.48 2.525 5.18 2.57 ;
      RECT 4.915 2.57 5.18 2.755 ;
      RECT 3.965 2.4 5.18 2.525 ;
      RECT 4.745 2.295 5.18 2.4 ;
      RECT 3.965 1.05 4.135 2.4 ;
      RECT 4.745 1.5 4.915 2.295 ;
      RECT 3.605 0.88 4.135 1.05 ;
      RECT 4.745 1.22 5.985 1.5 ;
      RECT 3.605 0.67 3.935 0.88 ;
      RECT 0 3.245 13.44 3.415 ;
      RECT 12.91 1.95 13.24 3.245 ;
      RECT 1 2.75 1.34 3.245 ;
      RECT 2.005 2.75 2.335 3.245 ;
      RECT 5.83 2.745 6.165 3.245 ;
      RECT 4.4 2.74 4.73 3.245 ;
      RECT 0.11 2.52 0.36 3.245 ;
      RECT 8.58 2.445 8.91 3.245 ;
      RECT 9.65 2.445 9.9 3.245 ;
      RECT 10.535 2.025 10.865 3.245 ;
      RECT 11.535 2.14 12.24 3.245 ;
      RECT 5.085 1.67 5.635 2.12 ;
      RECT 0.56 2.52 3.31 2.58 ;
      RECT 3.03 2.58 3.31 2.755 ;
      RECT 0.685 2.41 3.31 2.52 ;
      RECT 3.11 2.355 3.31 2.41 ;
      RECT 3.11 2.185 3.795 2.355 ;
      RECT 3.625 1.39 3.795 2.185 ;
      RECT 3.185 1.22 3.795 1.39 ;
      RECT 3.185 0.67 3.435 1.22 ;
      RECT 0.56 2.64 0.83 2.98 ;
      RECT 0.56 2.615 0.86 2.64 ;
      RECT 0.56 2.605 0.875 2.615 ;
      RECT 0.56 2.58 0.89 2.605 ;
      RECT 0.685 0.83 0.855 2.41 ;
      RECT 0.165 0.66 0.855 0.83 ;
      RECT 0.165 0.37 0.495 0.66 ;
      RECT 1.455 0.975 2.635 1.14 ;
      RECT 2.445 1.14 2.635 1.55 ;
      RECT 1.455 0.97 2.51 0.975 ;
      RECT 2.455 1.55 2.635 1.775 ;
      RECT 1.455 1.14 1.625 1.945 ;
      RECT 1.455 1.945 1.805 2.24 ;
      RECT 1.455 0.35 1.875 0.97 ;
      RECT 1.025 1.13 1.285 2.14 ;
      RECT 10.115 1.46 12.24 1.63 ;
      RECT 10.56 1.3 12.24 1.46 ;
      RECT 10.115 1.63 10.365 2.905 ;
      RECT 10.56 0.35 10.89 1.3 ;
      RECT 9.08 2.445 9.48 2.905 ;
      RECT 9.31 2.045 9.48 2.445 ;
      RECT 9.31 1.875 9.945 2.045 ;
      RECT 9.775 1.205 9.945 1.875 ;
      RECT 8.445 1.035 9.945 1.205 ;
      RECT 8.445 1.205 8.775 1.365 ;
      RECT 9.5 0.385 9.83 1.035 ;
      RECT 7.125 2.475 8.41 2.805 ;
      RECT 8.24 1.705 8.41 2.475 ;
      RECT 7.16 0.845 7.33 2.475 ;
      RECT 8.24 1.535 9.605 1.705 ;
      RECT 7.16 0.595 7.935 0.845 ;
      RECT 9.345 1.375 9.605 1.535 ;
      RECT 8.765 1.92 9.14 2.275 ;
      RECT 2.455 2.055 2.94 2.24 ;
      RECT 2.455 2.015 2.985 2.055 ;
      RECT 2.455 1.945 3.455 2.015 ;
      RECT 2.77 1.905 3.455 1.945 ;
      RECT 2.815 1.56 3.455 1.905 ;
      RECT 2.815 0.805 3.015 1.56 ;
      RECT 2.555 0.5 3.015 0.805 ;
      RECT 2.555 0.33 4.475 0.5 ;
      RECT 4.305 0.5 4.475 0.54 ;
      RECT 4.305 0.54 5.565 0.71 ;
      RECT 5.395 0.425 5.565 0.54 ;
      RECT 5.395 0.255 8.275 0.425 ;
      RECT 8.105 0.425 8.275 1.015 ;
      RECT 7.545 1.015 8.275 1.345 ;
      RECT 7.74 1.345 8.07 2.305 ;
      RECT 0 -0.085 13.44 0.085 ;
      RECT 13.005 0.085 13.335 1.1 ;
      RECT 1.065 0.085 1.235 0.83 ;
      RECT 2.055 0.085 2.385 0.8 ;
      RECT 4.895 0.085 5.225 0.37 ;
      RECT 8.625 0.085 8.955 0.845 ;
      RECT 10.115 0.085 10.39 1.13 ;
      RECT 11.12 0.085 11.41 1.13 ;
      RECT 12.08 0.085 12.405 0.71 ;
      RECT 6.155 1.94 6.615 2.235 ;
      RECT 6.155 1.05 6.325 1.94 ;
      RECT 4.305 0.88 6.99 1.05 ;
      RECT 4.305 1.05 4.57 2.105 ;
      RECT 5.735 0.72 6.99 0.88 ;
  END
END scs8ls_dfrtp_4

MACRO scs8ls_dfsbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.315 1.18 1.795 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475 1.01 0.805 2.02 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END D

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.12 1.18 10.435 2.98 ;
        RECT 10.12 1.13 10.315 1.18 ;
        RECT 9.985 0.35 10.315 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END QN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.555 1.82 11.885 2.98 ;
        RECT 11.715 1.05 11.885 1.82 ;
        RECT 11.555 0.35 11.885 1.05 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12 3.575 ;
    END
  END vpwr

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.375 1.595 8.545 1.735 ;
        RECT 5.375 1.735 5.665 1.78 ;
        RECT 8.255 1.735 8.545 1.78 ;
        RECT 5.375 1.55 5.665 1.595 ;
        RECT 8.255 1.55 8.545 1.595 ;
    END
    ANTENNAGATEAREA 0.252 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.205 LAYER met1 ;
  END SETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 5.435 1.58 5.605 1.75 ;
      RECT 8.315 1.58 8.485 1.75 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
    LAYER li1 ;
      RECT 9 2.56 9.33 2.98 ;
      RECT 9 2.39 9.735 2.56 ;
      RECT 9.565 1.01 9.735 2.39 ;
      RECT 7.77 0.84 9.735 1.01 ;
      RECT 7.77 1.01 8.1 1.88 ;
      RECT 8.925 0.415 9.255 0.84 ;
      RECT 0.975 1.89 1.455 2.02 ;
      RECT 0.975 1.72 2.355 1.89 ;
      RECT 2.025 1.3 2.355 1.72 ;
      RECT 0.975 0.35 1.435 1.01 ;
      RECT 0.975 1.01 1.145 1.72 ;
      RECT 8.285 1.18 8.67 1.78 ;
      RECT 0 3.245 12 3.415 ;
      RECT 11.05 1.995 11.38 3.245 ;
      RECT 9.56 2.73 9.91 3.245 ;
      RECT 8.07 2.65 8.24 3.245 ;
      RECT 0.565 2.59 0.895 3.245 ;
      RECT 1.575 2.53 1.905 3.245 ;
      RECT 4.045 2.505 4.44 3.245 ;
      RECT 5.71 2.465 6.05 3.245 ;
      RECT 0 -0.085 12 0.085 ;
      RECT 11.055 0.085 11.385 0.94 ;
      RECT 0.545 0.085 0.795 0.84 ;
      RECT 1.605 0.085 1.865 1.01 ;
      RECT 4.105 0.085 4.435 0.715 ;
      RECT 5.855 0.085 6.185 0.95 ;
      RECT 8.065 0.085 8.755 0.67 ;
      RECT 9.485 0.085 9.815 0.67 ;
      RECT 3.175 2.295 3.535 2.735 ;
      RECT 3.365 1.055 3.535 2.295 ;
      RECT 3.365 0.885 4.285 1.055 ;
      RECT 4.115 1.055 4.285 1.435 ;
      RECT 3.365 0.385 3.615 0.885 ;
      RECT 4.115 1.435 5.235 1.605 ;
      RECT 4.95 1.29 5.235 1.435 ;
      RECT 4.95 1.12 6.265 1.29 ;
      RECT 5.935 1.29 6.265 1.45 ;
      RECT 4.95 1.055 5.235 1.12 ;
      RECT 2.865 1.435 3.195 2.105 ;
      RECT 3.025 0.425 3.195 1.435 ;
      RECT 2.045 0.255 3.195 0.425 ;
      RECT 2.045 0.425 2.295 1.13 ;
      RECT 4.95 1.995 5.2 2.735 ;
      RECT 4.23 1.775 5.2 1.995 ;
      RECT 2.105 2.905 3.875 3.075 ;
      RECT 2.105 2.4 2.355 2.905 ;
      RECT 3.705 2.335 3.875 2.905 ;
      RECT 3.705 2.165 4.78 2.335 ;
      RECT 4.61 2.335 4.78 2.905 ;
      RECT 3.705 1.36 3.945 2.165 ;
      RECT 4.61 2.905 5.54 3.075 ;
      RECT 5.37 2.295 5.54 2.905 ;
      RECT 5.37 2.125 6.035 2.295 ;
      RECT 5.865 1.79 6.035 2.125 ;
      RECT 5.865 1.62 6.605 1.79 ;
      RECT 6.435 1.45 6.605 1.62 ;
      RECT 6.435 1.12 6.88 1.45 ;
      RECT 6.435 0.425 6.605 1.12 ;
      RECT 6.435 0.255 7.56 0.425 ;
      RECT 7.39 0.425 7.56 2.02 ;
      RECT 7.23 2.02 7.56 2.31 ;
      RECT 0.115 2.23 1.795 2.36 ;
      RECT 0.115 2.19 2.695 2.23 ;
      RECT 2.525 2.23 2.695 2.295 ;
      RECT 1.625 2.06 2.695 2.19 ;
      RECT 2.525 2.295 3.005 2.735 ;
      RECT 2.525 0.845 2.695 2.06 ;
      RECT 2.525 0.595 2.855 0.845 ;
      RECT 0.115 2.36 0.365 2.98 ;
      RECT 0.115 0.84 0.285 2.19 ;
      RECT 0.115 0.38 0.365 0.84 ;
      RECT 4.455 0.885 4.775 1.265 ;
      RECT 4.605 0.435 5.18 0.885 ;
      RECT 5.405 1.55 5.695 1.955 ;
      RECT 10.68 1.55 10.85 2.875 ;
      RECT 10.68 1.22 11.54 1.55 ;
      RECT 10.68 0.94 10.875 1.22 ;
      RECT 10.545 0.35 10.875 0.94 ;
      RECT 6.76 2.65 7.45 2.905 ;
      RECT 6.76 2.48 7.9 2.65 ;
      RECT 7.73 2.22 8.77 2.48 ;
      RECT 6.76 1.96 7.01 2.48 ;
      RECT 8.44 2.48 8.77 2.98 ;
      RECT 7.73 2.05 9.395 2.22 ;
      RECT 6.84 1.85 7.01 1.96 ;
      RECT 9.065 1.21 9.395 2.05 ;
      RECT 6.84 1.68 7.22 1.85 ;
      RECT 7.05 0.925 7.22 1.68 ;
      RECT 6.775 0.595 7.22 0.925 ;
  END
END scs8ls_dfsbp_1

MACRO scs8ls_dfsbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.085 0.35 12.425 1.13 ;
        RECT 12.255 1.13 12.425 1.82 ;
        RECT 12.065 1.82 12.425 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.175 0.35 10.435 1.82 ;
        RECT 10.13 1.82 10.435 2.97 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END QN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475 0.98 0.805 1.99 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.315 1.18 1.775 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END CLK

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12.96 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12.96 3.575 ;
    END
  END vpwr

  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.375 1.595 8.545 1.735 ;
        RECT 5.375 1.735 5.665 1.78 ;
        RECT 8.255 1.735 8.545 1.78 ;
        RECT 5.375 1.55 5.665 1.595 ;
        RECT 8.255 1.55 8.545 1.595 ;
    END
    ANTENNAGATEAREA 0.252 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.205 LAYER met1 ;
  END SETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 1.58 5.605 1.75 ;
      RECT 8.315 1.58 8.485 1.75 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
    LAYER li1 ;
      RECT 0.975 1.89 1.455 2.02 ;
      RECT 0.975 1.72 2.275 1.89 ;
      RECT 1.945 1.3 2.275 1.72 ;
      RECT 0.975 0.35 1.435 1.01 ;
      RECT 0.975 1.01 1.145 1.72 ;
      RECT 3.065 2.295 3.455 2.735 ;
      RECT 3.285 1.265 3.455 2.295 ;
      RECT 3.285 1.095 4.185 1.265 ;
      RECT 4.015 1.265 4.185 1.515 ;
      RECT 3.285 0.925 3.53 1.095 ;
      RECT 4.015 1.515 5.015 1.685 ;
      RECT 3.28 0.465 3.53 0.925 ;
      RECT 4.75 1.685 5.015 1.885 ;
      RECT 4.75 1.41 5.015 1.515 ;
      RECT 4.75 1.24 5.915 1.41 ;
      RECT 5.585 1.12 5.915 1.24 ;
      RECT 6.78 2.65 7.47 2.98 ;
      RECT 6.78 2.48 7.92 2.65 ;
      RECT 7.75 2.12 8.79 2.48 ;
      RECT 6.78 1.85 7.03 2.48 ;
      RECT 8.46 2.48 8.79 2.915 ;
      RECT 7.75 1.95 9.57 2.12 ;
      RECT 6.78 1.68 7.215 1.85 ;
      RECT 8.9 1.35 9.57 1.95 ;
      RECT 7.045 0.95 7.215 1.68 ;
      RECT 6.67 0.62 7.215 0.95 ;
      RECT 9.015 2.46 9.345 2.62 ;
      RECT 9.015 2.29 9.91 2.46 ;
      RECT 9.74 1.18 9.91 2.29 ;
      RECT 9.105 1.01 9.91 1.18 ;
      RECT 7.725 0.84 9.435 1.01 ;
      RECT 7.725 1.01 8.055 1.78 ;
      RECT 9.105 0.635 9.435 0.84 ;
      RECT 5.225 1.58 5.635 2.02 ;
      RECT 8.285 1.18 8.64 1.78 ;
      RECT 11.085 1.3 12.085 1.63 ;
      RECT 11.085 1.63 11.415 2.86 ;
      RECT 11.085 0.35 11.415 1.3 ;
      RECT 0 -0.085 12.96 0.085 ;
      RECT 12.595 0.085 12.845 1.13 ;
      RECT 10.605 0.085 10.855 1.13 ;
      RECT 11.585 0.085 11.915 1.03 ;
      RECT 0.545 0.085 0.795 0.81 ;
      RECT 1.605 0.085 1.865 1.01 ;
      RECT 3.99 0.085 4.24 0.845 ;
      RECT 5.34 0.085 6.16 0.68 ;
      RECT 8.1 0.085 8.845 0.67 ;
      RECT 9.665 0.085 9.995 0.84 ;
      RECT 0 3.245 12.96 3.415 ;
      RECT 12.595 1.82 12.845 3.245 ;
      RECT 10.605 1.82 10.86 3.245 ;
      RECT 11.615 1.82 11.865 3.245 ;
      RECT 4.02 2.735 4.35 3.245 ;
      RECT 8.09 2.65 8.26 3.245 ;
      RECT 9.63 2.63 9.96 3.245 ;
      RECT 0.565 2.53 0.895 3.245 ;
      RECT 1.575 2.53 1.905 3.245 ;
      RECT 5.7 2.53 6.07 3.245 ;
      RECT 4.355 1.015 4.58 1.345 ;
      RECT 4.41 0.35 4.88 1.015 ;
      RECT 2.785 1.435 3.115 2.105 ;
      RECT 2.94 0.425 3.11 1.435 ;
      RECT 2.045 0.255 3.11 0.425 ;
      RECT 2.045 0.425 2.215 1.13 ;
      RECT 4.86 2.295 5.19 2.735 ;
      RECT 4.86 2.225 5.03 2.295 ;
      RECT 4.14 2.055 5.03 2.225 ;
      RECT 4.14 1.855 4.47 2.055 ;
      RECT 2.105 2.905 3.845 3.075 ;
      RECT 3.625 2.565 3.845 2.905 ;
      RECT 2.105 2.4 2.275 2.905 ;
      RECT 3.625 2.395 4.69 2.565 ;
      RECT 4.52 2.565 4.69 2.905 ;
      RECT 3.625 1.435 3.845 2.395 ;
      RECT 4.52 2.905 5.53 3.075 ;
      RECT 5.36 2.36 5.53 2.905 ;
      RECT 5.36 2.19 6.5 2.36 ;
      RECT 6.33 1.45 6.5 2.19 ;
      RECT 6.33 1.12 6.875 1.45 ;
      RECT 6.33 0.45 6.5 1.12 ;
      RECT 6.33 0.28 7.555 0.45 ;
      RECT 7.385 0.45 7.555 2.02 ;
      RECT 7.25 2.02 7.58 2.31 ;
      RECT 0.115 2.23 1.795 2.36 ;
      RECT 0.115 2.19 2.615 2.23 ;
      RECT 2.445 2.23 2.615 2.295 ;
      RECT 1.625 2.06 2.615 2.19 ;
      RECT 2.445 2.295 2.865 2.735 ;
      RECT 2.445 0.925 2.615 2.06 ;
      RECT 2.445 0.595 2.77 0.925 ;
      RECT 0.115 2.36 0.365 2.98 ;
      RECT 0.115 0.81 0.285 2.19 ;
      RECT 0.115 0.35 0.365 0.81 ;
  END
END scs8ls_dfsbp_2

MACRO scs8ls_and3_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.45 3.23 1.78 ;
    END
    ANTENNAGATEAREA 0.444 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.325 4.335 1.78 ;
    END
    ANTENNAGATEAREA 0.444 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.615 1.45 5.285 1.78 ;
    END
    ANTENNAGATEAREA 0.444 ;
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.56 0.35 0.89 0.96 ;
        RECT 0.56 0.96 1.74 1.13 ;
        RECT 0.56 1.13 0.835 1.8 ;
        RECT 1.49 0.35 1.74 0.96 ;
        RECT 0.56 1.8 1.895 1.97 ;
        RECT 0.56 1.97 0.895 2.98 ;
        RECT 1.565 1.97 1.895 2.98 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 2.065 2.29 2.395 3.245 ;
      RECT 3.065 2.29 3.645 3.245 ;
      RECT 4.315 2.29 4.645 3.245 ;
      RECT 5.315 2.29 5.645 3.245 ;
      RECT 0.115 1.82 0.365 3.245 ;
      RECT 1.065 2.14 1.395 3.245 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 1.92 0.085 2.25 1.03 ;
      RECT 2.85 0.085 3.18 0.815 ;
      RECT 0.13 0.085 0.38 1.13 ;
      RECT 1.07 0.085 1.32 0.79 ;
      RECT 2.42 0.985 4.09 1.155 ;
      RECT 3.92 0.595 4.09 0.985 ;
      RECT 2.42 0.35 2.67 0.985 ;
      RECT 3.41 0.425 3.74 0.815 ;
      RECT 3.41 0.255 5.64 0.425 ;
      RECT 4.31 0.425 4.64 1.03 ;
      RECT 5.31 0.425 5.64 0.94 ;
      RECT 2.065 1.95 5.625 2.12 ;
      RECT 4.815 2.12 5.145 2.98 ;
      RECT 5.455 1.28 5.625 1.95 ;
      RECT 4.81 1.11 5.625 1.28 ;
      RECT 4.81 0.595 5.14 1.11 ;
      RECT 3.815 2.12 4.145 2.98 ;
      RECT 2.565 2.12 2.895 2.98 ;
      RECT 2.065 1.63 2.235 1.95 ;
      RECT 1.035 1.3 2.235 1.63 ;
    LAYER mcon ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_and3_4

MACRO scs8ls_and3b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005 1.39 2.335 1.78 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.39 2.875 1.78 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END C

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.11 0.57 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END AN

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.345 1.82 3.755 2.98 ;
        RECT 3.585 1.13 3.755 1.82 ;
        RECT 3.385 0.35 3.755 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.045 1.3 3.415 1.63 ;
      RECT 1.31 1.95 2.64 2.12 ;
      RECT 2.31 2.12 2.64 2.7 ;
      RECT 1.31 1.05 3.215 1.22 ;
      RECT 3.045 1.22 3.215 1.3 ;
      RECT 1.31 2.12 1.64 2.7 ;
      RECT 1.31 1.22 1.64 1.95 ;
      RECT 1.31 0.45 1.64 1.05 ;
      RECT 0.615 2.1 0.945 2.98 ;
      RECT 0.775 1.7 0.945 2.1 ;
      RECT 0.775 1.03 1.14 1.7 ;
      RECT 0.775 0.94 0.945 1.03 ;
      RECT 0.615 0.35 0.945 0.94 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 0.115 0.085 0.445 0.94 ;
      RECT 2.625 0.085 3.215 0.88 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 1.81 2.29 2.14 3.245 ;
      RECT 0.115 2.1 0.445 3.245 ;
      RECT 2.845 1.95 3.175 3.245 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_and3b_1

MACRO scs8ls_and3b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385 0.35 3.715 1.13 ;
        RECT 3.41 1.13 3.715 1.82 ;
        RECT 3.41 1.82 3.755 2.07 ;
    END
    ANTENNADIFFAREA 0.56 ;
  END X

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 0.44 2.45 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.69 1.35 3.235 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END C

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.26 0.55 1.93 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END AN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.42 2.24 4.215 2.41 ;
      RECT 4.045 1.63 4.215 2.24 ;
      RECT 3.885 1.3 4.215 1.63 ;
      RECT 2.42 2.41 2.75 2.86 ;
      RECT 2.42 2.12 2.75 2.24 ;
      RECT 1.4 1.95 2.75 2.12 ;
      RECT 1.4 2.12 1.73 2.86 ;
      RECT 1.4 0.35 1.755 1.95 ;
      RECT 0.115 2.27 0.4 2.98 ;
      RECT 0.115 2.1 1.07 2.27 ;
      RECT 0.9 1.855 1.07 2.1 ;
      RECT 0.9 1.09 1.23 1.855 ;
      RECT 0.115 0.92 1.23 1.09 ;
      RECT 0.115 0.42 0.375 0.92 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 3.895 0.085 4.145 1.13 ;
      RECT 2.815 0.085 3.145 1.13 ;
      RECT 0.545 0.085 0.875 0.75 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 2.96 2.58 3.29 3.245 ;
      RECT 3.875 2.58 4.205 3.245 ;
      RECT 0.57 2.44 0.9 3.245 ;
      RECT 1.9 2.29 2.23 3.245 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_and3b_2

MACRO scs8ls_and3b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.505 1.18 0.835 1.51 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END AN

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.35 3.56 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.55 6.595 1.8 ;
        RECT 4.57 1.8 6.595 1.97 ;
        RECT 4.57 1.97 4.9 2.98 ;
        RECT 5.57 1.97 5.9 2.98 ;
        RECT 5.935 1.13 6.105 1.8 ;
        RECT 4.965 0.96 6.105 1.13 ;
        RECT 4.965 0.35 5.215 0.96 ;
        RECT 5.925 0.35 6.105 0.96 ;
    END
    ANTENNADIFFAREA 1.1382 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 6.72 3.415 ;
      RECT 6.07 2.14 6.4 3.245 ;
      RECT 1.975 2.29 2.305 3.245 ;
      RECT 2.975 2.29 3.305 3.245 ;
      RECT 0.975 2.02 1.305 3.245 ;
      RECT 4.07 1.82 4.4 3.245 ;
      RECT 5.07 2.14 5.4 3.245 ;
      RECT 0 -0.085 6.72 0.085 ;
      RECT 6.275 0.085 6.605 1.13 ;
      RECT 0.615 0.085 0.875 1.01 ;
      RECT 3.525 0.085 3.855 0.84 ;
      RECT 4.465 0.085 4.795 1.13 ;
      RECT 5.395 0.085 5.725 0.79 ;
      RECT 2.035 0.72 2.365 1.15 ;
      RECT 2.035 0.47 3.295 0.72 ;
      RECT 2.035 0.425 2.365 0.47 ;
      RECT 1.175 0.255 2.365 0.425 ;
      RECT 1.175 0.425 1.505 1.15 ;
      RECT 2.535 1.01 4.285 1.18 ;
      RECT 2.535 0.89 2.865 1.01 ;
      RECT 4.035 0.45 4.285 1.01 ;
      RECT 0.475 1.85 0.805 2.86 ;
      RECT 0.115 1.68 1.305 1.85 ;
      RECT 1.135 1.65 1.305 1.68 ;
      RECT 1.135 1.32 1.525 1.65 ;
      RECT 0.115 1.01 0.285 1.68 ;
      RECT 0.115 0.35 0.445 1.01 ;
      RECT 3.73 1.46 5.765 1.63 ;
      RECT 4.755 1.3 5.765 1.46 ;
      RECT 1.475 1.95 3.9 2.12 ;
      RECT 3.535 2.12 3.9 2.86 ;
      RECT 3.73 1.63 3.9 1.95 ;
      RECT 2.475 2.12 2.805 2.86 ;
      RECT 1.475 2.12 1.805 2.86 ;
      RECT 1.475 1.82 1.865 1.95 ;
      RECT 1.695 1.15 1.865 1.82 ;
      RECT 1.685 0.595 1.865 1.15 ;
    LAYER mcon ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_and3b_4

MACRO scs8ls_and4_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.73 0.35 3.275 1.13 ;
        RECT 3.105 1.13 3.275 1.82 ;
        RECT 2.91 1.82 3.275 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 2.395 1.78 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END D

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.44 1.855 1.79 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985 0.44 1.315 1.805 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.12 0.815 1.79 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.57 1.32 2.935 1.65 ;
      RECT 0.085 2.13 2.205 2.145 ;
      RECT 1.875 2.145 2.205 2.98 ;
      RECT 0.085 1.975 2.74 2.13 ;
      RECT 1.875 1.96 2.74 1.975 ;
      RECT 2.57 1.65 2.74 1.96 ;
      RECT 0.615 2.145 0.945 2.98 ;
      RECT 0.085 0.355 0.77 0.95 ;
      RECT 0.085 0.95 0.255 1.975 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 0.115 2.315 0.445 3.245 ;
      RECT 1.115 2.315 1.705 3.245 ;
      RECT 2.41 2.3 2.74 3.245 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.22 0.085 2.55 1.03 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_and4_1

MACRO scs8ls_and4_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.79 0.77 3.235 1.13 ;
        RECT 2.835 1.13 3.235 2.15 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.3 0.445 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955 0.44 1.315 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.44 1.855 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.18 2.425 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.765 2.32 3.735 2.49 ;
      RECT 3.405 1.3 3.735 2.32 ;
      RECT 1.765 2.49 2.095 2.98 ;
      RECT 1.765 1.89 2.095 2.32 ;
      RECT 0.615 1.72 2.095 1.89 ;
      RECT 0.615 1.89 0.985 2.98 ;
      RECT 0.615 1.13 0.785 1.72 ;
      RECT 0.26 0.96 0.785 1.13 ;
      RECT 0.26 0.35 0.59 0.96 ;
      RECT 3.405 0.6 3.655 1.08 ;
      RECT 3.22 0.085 3.655 0.6 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 2.265 0.085 2.595 1.01 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 3.37 2.66 3.725 3.245 ;
      RECT 2.3 2.66 2.63 3.245 ;
      RECT 1.215 2.06 1.545 3.245 ;
      RECT 0.115 1.95 0.445 3.245 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_and4_2

MACRO scs8ls_and4_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.13 6.595 1.48 ;
        RECT 5.855 1.48 6.595 1.65 ;
        RECT 4.83 0.96 6.595 1.13 ;
        RECT 5.855 1.65 6.105 1.8 ;
        RECT 4.83 0.35 5.08 0.96 ;
        RECT 5.76 0.35 6.09 0.96 ;
        RECT 4.875 1.8 6.105 1.97 ;
        RECT 4.875 1.97 5.205 2.98 ;
        RECT 5.855 1.97 6.105 2.98 ;
    END
    ANTENNADIFFAREA 1.1646 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.06 1.45 1.39 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.45 0.55 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.98 1.345 4.365 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.93 1.47 3.26 1.8 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 4.535 1.3 5.685 1.63 ;
      RECT 2.43 1.97 4.705 2.12 ;
      RECT 2.43 2.12 4.145 2.14 ;
      RECT 3.815 1.95 4.705 1.97 ;
      RECT 3.815 2.14 4.145 2.98 ;
      RECT 4.535 1.63 4.705 1.95 ;
      RECT 1.56 2.24 1.73 2.98 ;
      RECT 0.565 1.95 1.73 2.24 ;
      RECT 1.56 1.77 1.73 1.95 ;
      RECT 1.56 1.6 2.76 1.77 ;
      RECT 0.72 1.005 1.33 1.255 ;
      RECT 2.43 1.77 2.76 1.97 ;
      RECT 2.43 2.14 2.76 2.98 ;
      RECT 0.72 1.255 0.89 1.95 ;
      RECT 0 -0.085 6.72 0.085 ;
      RECT 6.26 0.085 6.52 0.68 ;
      RECT 2.8 0.085 3.13 0.62 ;
      RECT 4.33 0.085 4.66 1.13 ;
      RECT 5.26 0.085 5.59 0.79 ;
      RECT 0 3.245 6.72 3.415 ;
      RECT 6.275 1.82 6.605 3.245 ;
      RECT 1.015 2.41 1.345 3.245 ;
      RECT 2.93 2.31 3.645 3.245 ;
      RECT 4.315 2.29 4.645 3.245 ;
      RECT 0.115 1.95 0.395 3.245 ;
      RECT 1.93 1.94 2.26 3.245 ;
      RECT 5.405 2.14 5.655 3.245 ;
      RECT 0.57 0.655 1.76 0.835 ;
      RECT 1.94 1.175 3.81 1.3 ;
      RECT 1.94 1.13 4.07 1.175 ;
      RECT 3.64 0.995 4.07 1.13 ;
      RECT 1.94 0.485 2.11 1.13 ;
      RECT 0.14 0.315 2.11 0.485 ;
      RECT 0.14 0.485 0.39 1.255 ;
      RECT 2.29 0.825 3.47 0.96 ;
      RECT 2.29 0.79 3.64 0.825 ;
      RECT 2.29 0.575 2.62 0.79 ;
      RECT 3.3 0.575 3.64 0.79 ;
    LAYER mcon ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_and4_4

MACRO scs8ls_and4b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.55 2.275 1.96 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 0.255 2.81 0.67 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985 1.55 3.315 1.88 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END D

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.19 0.595 1.86 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END AN

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.875 1.85 4.23 2.98 ;
        RECT 4.06 1.18 4.23 1.85 ;
        RECT 3.875 0.48 4.23 1.18 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.31 1.35 3.89 1.38 ;
      RECT 3.535 1.38 3.89 1.68 ;
      RECT 1.115 2.13 3.095 2.35 ;
      RECT 2.765 2.35 3.095 2.98 ;
      RECT 2.595 2.1 3.095 2.13 ;
      RECT 1.31 1.21 3.705 1.35 ;
      RECT 2.595 1.38 2.765 2.1 ;
      RECT 1.31 0.6 1.64 1.21 ;
      RECT 1.115 2.35 1.46 2.46 ;
      RECT 0.115 2.2 0.445 2.98 ;
      RECT 0.115 2.03 0.945 2.2 ;
      RECT 0.775 1.88 0.945 2.03 ;
      RECT 0.775 1.55 1.255 1.88 ;
      RECT 0.775 1.02 0.945 1.55 ;
      RECT 0.115 0.85 0.945 1.02 ;
      RECT 0.115 0.35 0.405 0.85 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 3.375 0.085 3.705 1.04 ;
      RECT 0.575 0.085 0.875 0.68 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 1.645 2.535 2.595 3.245 ;
      RECT 0.615 2.37 0.945 3.245 ;
      RECT 3.335 2.1 3.665 3.245 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_and4b_1

MACRO scs8ls_and4b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.35 3.405 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505 1.35 2.835 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965 1.35 2.295 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END D

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.3 0.455 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END AN

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055 1.82 1.44 2.2 ;
        RECT 1.055 1.13 1.225 1.82 ;
        RECT 1.055 0.35 1.385 1.13 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.61 1.95 3.645 2.2 ;
      RECT 1.61 0.96 4.07 1.13 ;
      RECT 3.74 0.35 4.07 0.96 ;
      RECT 1.61 1.63 1.78 1.95 ;
      RECT 1.395 1.3 1.78 1.63 ;
      RECT 1.61 1.13 1.78 1.3 ;
      RECT 0.115 2.37 3.985 2.54 ;
      RECT 3.815 1.68 3.985 2.37 ;
      RECT 3.615 1.35 3.985 1.68 ;
      RECT 0.115 2.54 0.445 2.7 ;
      RECT 0.115 1.95 0.795 2.37 ;
      RECT 0.625 1.13 0.795 1.95 ;
      RECT 0.115 0.96 0.795 1.13 ;
      RECT 0.115 0.54 0.445 0.96 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 1.555 0.085 2.165 0.79 ;
      RECT 0.625 0.085 0.875 0.79 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 0.65 2.71 0.98 3.245 ;
      RECT 1.645 2.71 1.975 3.245 ;
      RECT 2.74 2.71 3.07 3.245 ;
      RECT 3.85 2.71 4.205 3.245 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_and4b_2

MACRO scs8ls_and4b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 0.35 1.47 0.98 ;
        RECT 1.085 0.98 2.54 1.15 ;
        RECT 1.085 1.15 1.315 1.82 ;
        RECT 2.21 0.35 2.54 0.98 ;
        RECT 1.085 1.82 2.405 2.22 ;
    END
    ANTENNADIFFAREA 1.2096 ;
  END X

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845 1.47 7.18 1.8 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.915 1.35 3.245 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.47 5.155 1.8 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END D

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.19 0.835 1.55 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END AN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 5.655 0.765 5.905 0.96 ;
      RECT 5.655 0.595 6.955 0.765 ;
      RECT 6.625 0.765 6.955 0.935 ;
      RECT 3.46 1.18 5.475 1.3 ;
      RECT 3.3 1.13 5.475 1.18 ;
      RECT 3.3 0.605 3.63 1.13 ;
      RECT 5.305 0.425 5.475 1.13 ;
      RECT 5.305 0.255 7.495 0.425 ;
      RECT 7.165 0.425 7.495 0.96 ;
      RECT 3.81 0.79 5.125 0.96 ;
      RECT 3.81 0.63 4.105 0.79 ;
      RECT 4.795 0.605 5.125 0.79 ;
      RECT 2.575 1.97 6.88 2.22 ;
      RECT 5.65 1.94 6.08 1.97 ;
      RECT 5.91 1.3 6.08 1.94 ;
      RECT 5.91 1.13 6.335 1.3 ;
      RECT 6.08 0.935 6.335 1.13 ;
      RECT 2.575 1.95 3.515 1.97 ;
      RECT 2.575 1.65 2.745 1.95 ;
      RECT 1.485 1.32 2.745 1.65 ;
      RECT 0.085 2.39 7.52 2.56 ;
      RECT 7.35 1.3 7.52 2.39 ;
      RECT 6.505 1.13 7.52 1.3 ;
      RECT 6.505 1.3 6.675 1.47 ;
      RECT 6.25 1.47 6.675 1.8 ;
      RECT 0.085 2.56 0.445 2.86 ;
      RECT 0.085 1.82 0.445 2.39 ;
      RECT 0.085 1.02 0.255 1.82 ;
      RECT 0.085 0.45 0.405 1.02 ;
      RECT 0 -0.085 7.68 0.085 ;
      RECT 2.71 0.085 3.04 1.13 ;
      RECT 4.285 0.085 4.615 0.62 ;
      RECT 0.585 0.085 0.915 1.02 ;
      RECT 1.67 0.085 2 0.81 ;
      RECT 0 3.245 7.68 3.415 ;
      RECT 0.65 2.73 1.025 3.245 ;
      RECT 1.595 2.73 1.955 3.245 ;
      RECT 2.635 2.73 2.98 3.245 ;
      RECT 3.72 2.73 4.05 3.245 ;
      RECT 5.18 2.73 5.53 3.245 ;
      RECT 6.1 2.73 6.43 3.245 ;
      RECT 7 2.73 7.565 3.245 ;
    LAYER mcon ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
  END
END scs8ls_and4b_4

MACRO scs8ls_and4bb_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.3 0.4 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END AN

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.015 1.19 3.345 1.86 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END C

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.91 1.82 1.565 2.15 ;
        RECT 0.91 1.13 1.08 1.82 ;
        RECT 0.91 0.96 1.27 1.13 ;
        RECT 1.08 0.35 1.27 0.96 ;
    END
    ANTENNADIFFAREA 0.6925 ;
  END X

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.4 1.3 4.695 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END BN

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.515 1.19 3.89 1.86 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 4.315 2.12 4.645 2.98 ;
      RECT 4.06 1.95 4.645 2.12 ;
      RECT 4.06 1.02 4.685 1.03 ;
      RECT 2.555 0.85 4.685 1.02 ;
      RECT 4.355 0.44 4.685 0.85 ;
      RECT 4.06 1.03 4.23 1.95 ;
      RECT 2.555 1.02 2.845 1.79 ;
      RECT 2.215 2.03 3.625 2.2 ;
      RECT 3.295 2.2 3.625 2.98 ;
      RECT 2.295 2.2 2.625 2.98 ;
      RECT 2.215 1.03 2.385 2.03 ;
      RECT 1.44 0.86 2.385 1.03 ;
      RECT 1.44 1.03 1.61 1.3 ;
      RECT 1.82 0.35 2.385 0.86 ;
      RECT 1.25 1.3 1.61 1.63 ;
      RECT 0.115 2.32 2.045 2.49 ;
      RECT 1.78 1.29 2.045 2.32 ;
      RECT 0.115 2.49 0.445 2.7 ;
      RECT 0.115 1.95 0.74 2.32 ;
      RECT 0.57 1.13 0.74 1.95 ;
      RECT 0.115 0.96 0.74 1.13 ;
      RECT 0.115 0.35 0.365 0.96 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 0.65 2.66 0.98 3.245 ;
      RECT 1.795 2.66 2.125 3.245 ;
      RECT 2.795 2.37 3.125 3.245 ;
      RECT 3.815 2.29 4.145 3.245 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 3.72 0.085 4.11 0.68 ;
      RECT 0.545 0.085 0.875 0.79 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_and4bb_1

MACRO scs8ls_and4bb_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.31 1.42 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.42 3.255 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END D

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.45 0.55 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END AN

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.825 1.18 5.155 1.59 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END BN

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.835 1.84 4.195 2.98 ;
        RECT 4.025 1.17 4.195 1.84 ;
        RECT 3.815 0.92 4.195 1.17 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 5.28 3.415 ;
      RECT 4.365 2.1 4.615 3.245 ;
      RECT 0.78 2.29 1.11 3.245 ;
      RECT 2.065 2.29 2.395 3.245 ;
      RECT 3.2 2.29 3.53 3.245 ;
      RECT 0.21 2.12 0.54 2.82 ;
      RECT 0.21 1.95 0.935 2.12 ;
      RECT 0.765 1.67 0.935 1.95 ;
      RECT 0.765 1.34 1.26 1.67 ;
      RECT 0.765 1.28 0.935 1.34 ;
      RECT 0.115 1.11 0.935 1.28 ;
      RECT 0.115 0.35 0.365 1.11 ;
      RECT 4.82 1.93 5.165 2.7 ;
      RECT 4.365 1.76 5.165 1.93 ;
      RECT 3.475 0.58 5.165 0.75 ;
      RECT 4.835 0.75 5.165 1.01 ;
      RECT 4.365 0.75 4.535 1.76 ;
      RECT 3.475 0.75 3.645 1 ;
      RECT 1.77 1 3.645 1.17 ;
      RECT 1.77 1.17 2.1 1.59 ;
      RECT 3.495 1.34 3.855 1.67 ;
      RECT 1.43 1.95 3.665 2.12 ;
      RECT 2.61 2.12 2.94 2.98 ;
      RECT 3.495 1.67 3.665 1.95 ;
      RECT 1.43 2.12 1.76 2.98 ;
      RECT 1.43 1.94 1.76 1.95 ;
      RECT 1.43 1.17 1.6 1.94 ;
      RECT 1.105 0.39 1.6 1.17 ;
      RECT 0 -0.085 5.28 0.085 ;
      RECT 4.325 0.085 4.655 0.41 ;
      RECT 0.545 0.085 0.875 0.94 ;
      RECT 2.975 0.085 3.305 0.83 ;
    LAYER mcon ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_and4bb_2

MACRO scs8ls_and4bb_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.24 0.77 8.995 0.98 ;
        RECT 7.24 0.98 8.995 1.15 ;
        RECT 8.765 1.15 8.995 1.82 ;
        RECT 7.24 0.35 7.57 0.98 ;
        RECT 7.405 1.82 8.995 2.15 ;
        RECT 7.405 2.15 7.575 2.98 ;
    END
    ANTENNADIFFAREA 1.116 ;
  END X

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.965 1.45 6.115 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END C

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.35 6.875 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END D

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.45 1.335 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END AN

  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.45 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END BN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.045 0.585 1.53 0.94 ;
      RECT 1.045 0.255 1.69 0.585 ;
      RECT 2.04 1.095 2.37 1.28 ;
      RECT 2.2 0.925 2.37 1.095 ;
      RECT 2.2 0.755 3.22 0.925 ;
      RECT 3.05 0.925 3.22 1.255 ;
      RECT 3.05 1.255 4.16 1.425 ;
      RECT 3.83 1.095 4.16 1.255 ;
      RECT 3.4 0.925 3.65 1.085 ;
      RECT 3.4 0.755 5.22 0.925 ;
      RECT 4.89 0.925 5.22 0.94 ;
      RECT 4.89 0.665 5.22 0.755 ;
      RECT 4.39 1.28 4.72 1.345 ;
      RECT 4.39 1.18 5.65 1.28 ;
      RECT 4.39 1.11 6.56 1.18 ;
      RECT 4.39 1.095 4.72 1.11 ;
      RECT 5.4 1.01 6.56 1.11 ;
      RECT 5.4 0.665 5.65 1.01 ;
      RECT 6.31 0.45 6.56 1.01 ;
      RECT 1.115 2.46 1.445 2.98 ;
      RECT 1.115 2.29 2.26 2.46 ;
      RECT 1.93 1.45 2.26 2.29 ;
      RECT 7.065 1.32 8.565 1.65 ;
      RECT 4.465 1.95 7.235 2.12 ;
      RECT 6.335 2.12 6.665 2.86 ;
      RECT 7.065 1.65 7.235 1.95 ;
      RECT 4.465 2.12 4.795 2.96 ;
      RECT 4.465 1.765 4.795 1.95 ;
      RECT 2.43 1.595 4.795 1.765 ;
      RECT 2.43 1.765 2.76 2.96 ;
      RECT 3.465 1.765 3.795 2.96 ;
      RECT 2.54 1.36 2.76 1.595 ;
      RECT 2.54 1.095 2.87 1.36 ;
      RECT 0.115 1.95 1.675 2.12 ;
      RECT 1.505 1.28 1.675 1.95 ;
      RECT 0.115 1.11 1.87 1.28 ;
      RECT 1.7 0.925 1.87 1.11 ;
      RECT 1.7 0.755 2.03 0.925 ;
      RECT 1.86 0.585 2.03 0.755 ;
      RECT 1.86 0.255 3.605 0.585 ;
      RECT 0.115 2.12 0.445 2.98 ;
      RECT 0.115 0.35 0.365 1.11 ;
      RECT 0 -0.085 9.12 0.085 ;
      RECT 8.67 0.085 9.005 0.6 ;
      RECT 0.545 0.085 0.875 0.94 ;
      RECT 5.88 0.085 6.13 0.84 ;
      RECT 6.74 0.085 7.07 1.13 ;
      RECT 7.74 0.085 8.07 0.81 ;
      RECT 0 3.245 9.12 3.415 ;
      RECT 7.775 2.32 8.105 3.245 ;
      RECT 8.675 2.32 9.005 3.245 ;
      RECT 1.89 2.63 2.225 3.245 ;
      RECT 0.615 2.29 0.945 3.245 ;
      RECT 4.965 2.29 6.165 3.245 ;
      RECT 6.875 2.29 7.205 3.245 ;
      RECT 2.965 1.935 3.295 3.245 ;
      RECT 3.965 1.935 4.295 3.245 ;
    LAYER mcon ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
  END
END scs8ls_and4bb_4

MACRO scs8ls_buf_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.47 1.82 1.83 2.98 ;
        RECT 1.66 1.13 1.83 1.82 ;
        RECT 1.475 0.35 1.83 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.45 0.91 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.13 1.3 1.49 1.63 ;
      RECT 0.47 2.12 0.8 2.98 ;
      RECT 0.47 1.95 1.3 2.12 ;
      RECT 1.13 1.63 1.3 1.95 ;
      RECT 1.13 1.28 1.3 1.3 ;
      RECT 0.115 1.11 1.3 1.28 ;
      RECT 0.115 0.8 0.795 1.11 ;
      RECT 0 -0.085 1.92 0.085 ;
      RECT 0.975 0.085 1.305 0.94 ;
      RECT 0 3.245 1.92 3.415 ;
      RECT 0.97 2.29 1.3 3.245 ;
    LAYER mcon ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_buf_1

MACRO scs8ls_buf_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.775 1.35 10.435 1.78 ;
    END
    ANTENNAGATEAREA 1.674 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
    END
  END vpwr

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.575 1.92 7.255 2.15 ;
    END
    ANTENNADIFFAREA 4.3456 ;
  END X

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 0.985 1.55 7.65 1.78 ;
    LAYER li1 ;
      RECT 0.13 0.085 0.38 1.13 ;
      RECT 0 -0.085 10.56 0.085 ;
      RECT 0.99 0.085 1.285 1.13 ;
      RECT 1.895 0.085 2.1 1.13 ;
      RECT 2.79 0.085 2.96 1.015 ;
      RECT 3.65 0.085 3.82 1.13 ;
      RECT 4.555 0.085 4.83 1.13 ;
      RECT 5.5 0.085 5.83 1.035 ;
      RECT 6.5 0.085 6.83 1.13 ;
      RECT 7.43 0.085 7.76 0.84 ;
      RECT 8.29 0.085 8.62 0.84 ;
      RECT 9.15 0.085 9.48 0.84 ;
      RECT 10.115 0.085 10.445 1.13 ;
      RECT 0 3.245 10.56 3.415 ;
      RECT 7.445 2.29 7.695 3.245 ;
      RECT 8.395 2.29 8.565 3.245 ;
      RECT 9.295 2.29 9.465 3.245 ;
      RECT 1.095 1.965 1.265 3.245 ;
      RECT 1.965 1.965 2.215 3.245 ;
      RECT 2.945 1.965 3.115 3.245 ;
      RECT 3.845 1.965 4.015 3.245 ;
      RECT 4.745 1.965 4.915 3.245 ;
      RECT 5.645 1.965 5.815 3.245 ;
      RECT 6.545 1.965 6.715 3.245 ;
      RECT 10.195 1.95 10.445 3.245 ;
      RECT 0.115 1.82 0.365 3.245 ;
      RECT 7.865 2.12 8.195 2.98 ;
      RECT 7.42 1.95 9.995 2.12 ;
      RECT 8.765 2.12 9.095 2.98 ;
      RECT 9.665 2.12 9.995 2.98 ;
      RECT 7.42 1.01 9.945 1.18 ;
      RECT 7.94 0.35 8.11 1.01 ;
      RECT 8.8 0.35 8.97 1.01 ;
      RECT 9.695 0.35 9.945 1.01 ;
      RECT 7.42 1.18 7.59 1.95 ;
      RECT 6.98 1.25 7.245 2.98 ;
      RECT 7 0.35 7.25 1.25 ;
      RECT 6.06 1.13 6.33 2.98 ;
      RECT 6 0.35 6.33 1.13 ;
      RECT 5.115 1.375 5.41 2.98 ;
      RECT 5.035 1.205 5.41 1.375 ;
      RECT 5.035 0.35 5.33 1.205 ;
      RECT 4.215 1.9 4.545 2.98 ;
      RECT 4.215 1.13 4.385 1.9 ;
      RECT 4 0.35 4.385 1.13 ;
      RECT 0.985 1.3 1.295 1.78 ;
      RECT 1.89 1.3 2.175 1.78 ;
      RECT 2.845 1.3 3.14 1.78 ;
      RECT 3.735 1.655 4.045 1.78 ;
      RECT 3.655 1.3 4.045 1.655 ;
      RECT 4.675 1.73 4.865 1.78 ;
      RECT 4.555 1.3 4.865 1.73 ;
      RECT 5.58 1.3 5.89 1.78 ;
      RECT 6.5 1.3 6.81 1.78 ;
      RECT 3.31 1.82 3.565 2.98 ;
      RECT 3.31 1.13 3.48 1.82 ;
      RECT 3.22 0.35 3.48 1.13 ;
      RECT 2.415 1.355 2.675 2.98 ;
      RECT 2.345 1.185 2.675 1.355 ;
      RECT 2.345 0.35 2.61 1.185 ;
      RECT 1.465 0.35 1.72 2.98 ;
      RECT 0.56 0.35 0.815 2.98 ;
    LAYER mcon ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 0.635 1.95 0.805 2.12 ;
      RECT 1.515 1.95 1.685 2.12 ;
      RECT 2.47 1.95 2.64 2.12 ;
      RECT 3.36 1.95 3.53 2.12 ;
      RECT 4.3 1.95 4.47 2.12 ;
      RECT 5.195 1.95 5.365 2.12 ;
      RECT 6.095 1.95 6.265 2.12 ;
      RECT 7.025 1.95 7.195 2.12 ;
      RECT 6.565 1.58 6.735 1.75 ;
      RECT 5.65 1.58 5.82 1.75 ;
      RECT 4.68 1.58 4.85 1.75 ;
      RECT 3.8 1.58 3.97 1.75 ;
      RECT 2.91 1.58 3.08 1.75 ;
      RECT 1.95 1.58 2.12 1.75 ;
      RECT 1.055 1.58 1.225 1.75 ;
      RECT 7.42 1.58 7.59 1.75 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
  END
END scs8ls_buf_16

MACRO scs8ls_buf_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 1.18 1.315 2.15 ;
        RECT 0.945 0.35 1.275 1.18 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.825 1.35 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 2.4 3.415 ;
      RECT 1.395 2.66 1.725 3.245 ;
      RECT 0.115 2.735 0.825 3.245 ;
      RECT 0.115 1.82 0.42 2.735 ;
      RECT 1.93 2.49 2.285 2.88 ;
      RECT 0.605 2.32 2.285 2.49 ;
      RECT 1.93 1.95 2.285 2.32 ;
      RECT 1.485 1.01 2.285 1.18 ;
      RECT 1.955 0.45 2.285 1.01 ;
      RECT 1.485 1.18 1.655 2.32 ;
      RECT 0.605 1.63 0.775 2.32 ;
      RECT 0.105 1.3 0.775 1.63 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 1.445 0.085 1.775 0.84 ;
      RECT 0.515 0.085 0.765 1.13 ;
    LAYER mcon ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_buf_2

MACRO scs8ls_buf_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.18 0.835 1.41 ;
        RECT 0.66 1.41 0.835 1.8 ;
        RECT 0.615 1.13 0.835 1.18 ;
        RECT 0.66 1.8 1.73 1.97 ;
        RECT 0.615 0.96 1.945 1.13 ;
        RECT 0.66 1.97 0.835 2.98 ;
        RECT 1.56 1.97 1.73 2.98 ;
        RECT 0.615 0.35 0.945 0.96 ;
        RECT 1.615 0.35 1.945 0.96 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.35 2.905 1.78 ;
    END
    ANTENNAGATEAREA 0.363 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.465 1.95 3.245 2.2 ;
      RECT 3.075 1.13 3.245 1.95 ;
      RECT 2.115 0.96 3.245 1.13 ;
      RECT 2.915 0.35 3.245 0.96 ;
      RECT 2.115 1.13 2.285 1.3 ;
      RECT 1.06 1.3 2.285 1.63 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.915 2.37 3.245 3.245 ;
      RECT 1.93 1.82 2.26 3.245 ;
      RECT 0.13 1.82 0.46 3.245 ;
      RECT 1.03 2.14 1.36 3.245 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.115 0.085 2.745 0.68 ;
      RECT 0.115 0.085 0.445 1.01 ;
      RECT 1.115 0.085 1.445 0.79 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_buf_4

MACRO scs8ls_buf_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.43 1.78 ;
    END
    ANTENNAGATEAREA 0.837 ;
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.82 1.97 5.155 2.98 ;
        RECT 1.97 1.8 5.155 1.97 ;
        RECT 1.97 1.97 2.3 2.98 ;
        RECT 2.92 1.97 3.25 2.98 ;
        RECT 3.87 1.97 4.2 2.98 ;
        RECT 4.975 1.13 5.145 1.8 ;
        RECT 1.96 0.96 5.145 1.13 ;
        RECT 1.96 0.35 2.13 0.96 ;
        RECT 2.81 0.35 3.14 0.96 ;
        RECT 3.81 0.35 4.14 0.96 ;
        RECT 4.81 0.35 5.145 0.96 ;
    END
    ANTENNADIFFAREA 2.2493 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.6 1.3 4.805 1.63 ;
      RECT 0.12 2.12 0.45 2.98 ;
      RECT 0.12 1.95 1.77 2.12 ;
      RECT 1.02 2.12 1.35 2.98 ;
      RECT 1.6 1.63 1.77 1.95 ;
      RECT 1.6 1.18 1.77 1.3 ;
      RECT 0.115 1.01 1.77 1.18 ;
      RECT 0.115 0.35 0.365 1.01 ;
      RECT 1.1 0.35 1.27 1.01 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 5.35 1.82 5.6 3.245 ;
      RECT 0.65 2.29 0.82 3.245 ;
      RECT 1.55 2.29 1.8 3.245 ;
      RECT 2.5 2.14 2.75 3.245 ;
      RECT 3.45 2.14 3.7 3.245 ;
      RECT 4.4 2.14 4.65 3.245 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 5.315 0.085 5.645 1.13 ;
      RECT 0.545 0.085 0.875 0.84 ;
      RECT 1.45 0.085 1.78 0.84 ;
      RECT 2.31 0.085 2.64 0.79 ;
      RECT 3.31 0.085 3.64 0.79 ;
      RECT 4.31 0.085 4.64 0.79 ;
    LAYER mcon ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_buf_8

MACRO scs8ls_bufbuf_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.3 0.505 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12.96 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12.96 3.575 ;
    END
  END vpwr

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.7 1.92 12.38 2.15 ;
    END
    ANTENNADIFFAREA 4.4016 ;
  END X

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 7 1.58 7.17 1.75 ;
      RECT 6.125 1.58 6.295 1.75 ;
      RECT 5.18 1.58 5.35 1.75 ;
      RECT 11.6 1.58 11.77 1.75 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.76 1.95 5.93 2.12 ;
      RECT 6.675 1.95 6.845 2.12 ;
      RECT 7.595 1.95 7.765 2.12 ;
      RECT 8.485 1.95 8.655 2.12 ;
      RECT 9.405 1.95 9.575 2.12 ;
      RECT 10.295 1.95 10.465 2.12 ;
      RECT 11.195 1.95 11.365 2.12 ;
      RECT 12.115 1.95 12.285 2.12 ;
      RECT 10.675 1.58 10.845 1.75 ;
      RECT 9.73 1.58 9.9 1.75 ;
      RECT 8.82 1.58 8.99 1.75 ;
      RECT 7.9 1.58 8.07 1.75 ;
    LAYER met1 ;
      RECT 5.11 1.55 11.83 1.78 ;
    LAYER li1 ;
      RECT 0 3.245 12.96 3.415 ;
      RECT 0.645 2.29 0.815 3.245 ;
      RECT 3.47 2.16 3.64 3.245 ;
      RECT 4.37 2.16 4.54 3.245 ;
      RECT 1.545 2.14 1.715 3.245 ;
      RECT 5.28 1.925 5.45 3.245 ;
      RECT 6.16 1.925 6.41 3.245 ;
      RECT 7.14 1.925 7.31 3.245 ;
      RECT 8.04 1.925 8.21 3.245 ;
      RECT 8.94 1.925 9.11 3.245 ;
      RECT 9.84 1.925 10.01 3.245 ;
      RECT 10.74 1.925 10.91 3.245 ;
      RECT 11.64 1.925 11.89 3.245 ;
      RECT 2.49 1.82 2.74 3.245 ;
      RECT 12.59 1.82 12.84 3.245 ;
      RECT 0.56 0.085 0.89 0.79 ;
      RECT 0 -0.085 12.96 0.085 ;
      RECT 1.42 0.085 1.67 0.79 ;
      RECT 2.415 0.085 2.745 1.13 ;
      RECT 3.345 0.085 3.675 0.81 ;
      RECT 4.275 0.085 4.605 0.81 ;
      RECT 5.275 0.085 5.455 1.13 ;
      RECT 6.065 0.085 6.315 1.13 ;
      RECT 6.96 0.085 7.175 1.13 ;
      RECT 7.85 0.085 8.115 1.13 ;
      RECT 8.75 0.085 9.045 1.13 ;
      RECT 9.665 0.085 9.975 1.13 ;
      RECT 10.575 0.085 10.905 1.13 ;
      RECT 11.505 0.085 11.835 1.13 ;
      RECT 12.515 0.085 12.845 1.13 ;
      RECT 6.055 1.32 6.365 1.75 ;
      RECT 6.95 1.32 7.215 1.75 ;
      RECT 7.85 1.32 8.115 1.75 ;
      RECT 8.75 1.32 9.045 1.75 ;
      RECT 9.65 1.32 9.975 1.75 ;
      RECT 10.565 1.32 10.94 1.75 ;
      RECT 11.495 1.32 11.89 1.75 ;
      RECT 5.66 1.92 5.99 2.98 ;
      RECT 5.66 1.9 5.885 1.92 ;
      RECT 5.635 0.35 5.885 1.9 ;
      RECT 2.94 1.99 3.27 2.98 ;
      RECT 2.94 1.82 5.08 1.99 ;
      RECT 3.84 1.99 4.17 2.98 ;
      RECT 4.75 1.99 5.08 2.98 ;
      RECT 4.845 1.755 5.08 1.82 ;
      RECT 4.845 1.32 5.405 1.755 ;
      RECT 4.845 1.15 5.105 1.32 ;
      RECT 2.915 0.98 5.105 1.15 ;
      RECT 2.915 0.35 3.165 0.98 ;
      RECT 3.845 0.35 4.095 0.98 ;
      RECT 4.775 0.35 5.025 0.98 ;
      RECT 1.015 1.97 1.345 2.98 ;
      RECT 1.015 1.8 2.245 1.97 ;
      RECT 1.915 1.97 2.245 2.98 ;
      RECT 2.045 1.65 2.245 1.8 ;
      RECT 2.045 1.32 4.48 1.65 ;
      RECT 2.045 1.13 2.215 1.32 ;
      RECT 1.07 0.96 2.215 1.13 ;
      RECT 1.07 0.35 1.24 0.96 ;
      RECT 1.855 0.35 2.215 0.96 ;
      RECT 0.115 2.12 0.445 2.98 ;
      RECT 0.115 1.95 0.845 2.12 ;
      RECT 0.675 1.63 0.845 1.95 ;
      RECT 0.675 1.3 1.875 1.63 ;
      RECT 0.675 1.13 0.845 1.3 ;
      RECT 0.13 0.96 0.845 1.13 ;
      RECT 0.13 0.35 0.38 0.96 ;
      RECT 12.06 2.02 12.39 2.98 ;
      RECT 12.06 1.15 12.345 2.02 ;
      RECT 12.015 0.35 12.345 1.15 ;
      RECT 11.11 1.92 11.44 2.98 ;
      RECT 11.11 0.35 11.325 1.92 ;
      RECT 10.21 1.92 10.54 2.98 ;
      RECT 10.21 1.65 10.395 1.92 ;
      RECT 10.145 0.35 10.395 1.65 ;
      RECT 9.31 1.92 9.64 2.98 ;
      RECT 9.31 1.65 9.48 1.92 ;
      RECT 9.215 0.35 9.48 1.65 ;
      RECT 8.41 1.92 8.74 2.98 ;
      RECT 8.41 1.65 8.58 1.92 ;
      RECT 8.285 0.35 8.58 1.65 ;
      RECT 7.51 1.92 7.84 2.98 ;
      RECT 7.51 1.65 7.68 1.92 ;
      RECT 7.385 0.35 7.68 1.65 ;
      RECT 6.61 1.92 6.94 2.98 ;
      RECT 6.61 1.65 6.78 1.92 ;
      RECT 6.535 0.35 6.78 1.65 ;
  END
END scs8ls_bufbuf_16

MACRO scs8ls_bufbuf_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.255 1.27 7.075 1.78 ;
        RECT 6.255 1.78 6.555 1.8 ;
        RECT 6.255 1.13 6.585 1.27 ;
        RECT 3.565 1.8 6.555 1.97 ;
        RECT 3.475 0.88 6.585 1.13 ;
        RECT 3.565 1.97 3.83 2.98 ;
        RECT 4.495 1.97 4.745 2.98 ;
        RECT 5.385 1.97 5.655 2.98 ;
        RECT 6.285 1.97 6.555 2.98 ;
        RECT 3.475 0.35 3.805 0.88 ;
        RECT 6.255 0.35 6.585 0.88 ;
    END
    ANTENNADIFFAREA 2.2732 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 0.57 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 7.2 0.085 ;
      RECT 6.755 0.085 7.085 1.1 ;
      RECT 0.625 0.085 0.955 0.84 ;
      RECT 2.115 0.085 2.445 0.71 ;
      RECT 2.975 0.085 3.305 0.71 ;
      RECT 3.975 0.085 4.305 0.71 ;
      RECT 4.835 0.085 5.165 0.71 ;
      RECT 5.755 0.085 6.085 0.71 ;
      RECT 0 3.245 7.2 3.415 ;
      RECT 6.735 1.95 7.04 3.245 ;
      RECT 0.565 2.37 0.92 3.245 ;
      RECT 2.15 2.16 2.38 3.245 ;
      RECT 3.05 1.82 3.38 3.245 ;
      RECT 4.035 2.14 4.29 3.245 ;
      RECT 4.93 2.14 5.205 3.245 ;
      RECT 5.835 2.14 6.105 3.245 ;
      RECT 0.115 2.2 0.38 2.7 ;
      RECT 0.115 1.95 0.92 2.2 ;
      RECT 0.75 1.63 0.92 1.95 ;
      RECT 0.75 1.3 1.14 1.63 ;
      RECT 0.75 1.18 0.92 1.3 ;
      RECT 0.115 1.01 0.92 1.18 ;
      RECT 0.115 0.54 0.445 1.01 ;
      RECT 2.67 1.3 6.02 1.63 ;
      RECT 1.65 1.99 1.98 2.98 ;
      RECT 1.65 1.82 2.88 1.99 ;
      RECT 2.55 1.99 2.88 2.98 ;
      RECT 2.67 1.63 2.88 1.82 ;
      RECT 2.67 1.13 3.125 1.3 ;
      RECT 1.685 0.88 3.125 1.13 ;
      RECT 1.685 0.35 1.935 0.88 ;
      RECT 1.09 1.82 1.48 2.98 ;
      RECT 1.31 1.63 1.48 1.82 ;
      RECT 1.31 1.3 2.5 1.63 ;
      RECT 1.31 1.13 1.48 1.3 ;
      RECT 1.125 0.35 1.48 1.13 ;
    LAYER mcon ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_bufbuf_8

MACRO scs8ls_bufinv_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.43 1.78 ;
    END
    ANTENNAGATEAREA 0.837 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 12 3.575 ;
    END
  END vpwr

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.66 1.92 11.4 2.15 ;
    END
    ANTENNADIFFAREA 4.3904 ;
  END Y

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.92 1.58 7.09 1.75 ;
      RECT 5.98 1.58 6.15 1.75 ;
      RECT 5.09 1.58 5.26 1.75 ;
      RECT 4.225 1.58 4.395 1.75 ;
      RECT 10.625 1.58 10.795 1.75 ;
      RECT 11.17 1.95 11.34 2.12 ;
      RECT 10.22 1.95 10.39 2.12 ;
      RECT 9.27 1.95 9.44 2.12 ;
      RECT 8.32 1.95 8.49 2.12 ;
      RECT 7.42 1.95 7.59 2.12 ;
      RECT 6.52 1.95 6.69 2.12 ;
      RECT 5.62 1.95 5.79 2.12 ;
      RECT 4.73 1.95 4.9 2.12 ;
      RECT 9.69 1.58 9.86 1.75 ;
      RECT 8.765 1.58 8.935 1.75 ;
      RECT 7.835 1.58 8.005 1.75 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
    LAYER met1 ;
      RECT 4.155 1.55 10.855 1.78 ;
    LAYER li1 ;
      RECT 5.035 1.3 5.305 1.75 ;
      RECT 5.9 1.3 6.23 1.75 ;
      RECT 6.84 1.3 7.17 1.75 ;
      RECT 7.76 1.3 8.09 1.75 ;
      RECT 8.685 1.3 9.015 1.75 ;
      RECT 9.615 1.3 9.945 1.75 ;
      RECT 10.545 1.3 10.875 1.75 ;
      RECT 0.12 2.12 0.45 2.98 ;
      RECT 0.12 1.95 1.77 2.12 ;
      RECT 1.02 2.12 1.35 2.98 ;
      RECT 1.6 1.63 1.77 1.95 ;
      RECT 1.6 1.3 3.46 1.63 ;
      RECT 1.6 1.18 1.77 1.3 ;
      RECT 0.115 1.01 1.77 1.18 ;
      RECT 0.115 0.35 0.365 1.01 ;
      RECT 1.115 0.35 1.285 1.01 ;
      RECT 1.94 1.97 2.27 2.98 ;
      RECT 1.94 1.8 4.07 1.97 ;
      RECT 2.84 1.97 3.17 2.98 ;
      RECT 3.74 1.97 4.07 2.98 ;
      RECT 3.74 1.75 4.07 1.8 ;
      RECT 3.74 1.3 4.435 1.75 ;
      RECT 3.685 1.13 3.935 1.3 ;
      RECT 1.975 0.96 3.935 1.13 ;
      RECT 1.975 0.35 2.145 0.96 ;
      RECT 2.755 0.35 3.005 0.96 ;
      RECT 3.685 0.35 3.935 0.96 ;
      RECT 0 3.245 12 3.415 ;
      RECT 0.65 2.29 0.82 3.245 ;
      RECT 1.55 2.29 1.72 3.245 ;
      RECT 2.47 2.14 2.64 3.245 ;
      RECT 3.37 2.14 3.54 3.245 ;
      RECT 4.27 1.92 4.44 3.245 ;
      RECT 5.17 1.92 5.34 3.245 ;
      RECT 6.07 1.92 6.24 3.245 ;
      RECT 6.97 1.92 7.14 3.245 ;
      RECT 7.87 1.92 8.04 3.245 ;
      RECT 8.77 1.92 8.995 3.245 ;
      RECT 9.72 1.92 9.955 3.245 ;
      RECT 10.67 1.92 10.885 3.245 ;
      RECT 11.62 1.82 11.87 3.245 ;
      RECT 11.09 2.02 11.42 2.98 ;
      RECT 11.055 1.79 11.42 2.02 ;
      RECT 11.055 0.35 11.385 1.79 ;
      RECT 0.545 0.085 0.875 0.84 ;
      RECT 0 -0.085 12 0.085 ;
      RECT 1.465 0.085 1.795 0.84 ;
      RECT 2.325 0.085 2.575 0.79 ;
      RECT 3.185 0.085 3.515 0.79 ;
      RECT 4.115 0.085 4.445 1.13 ;
      RECT 5.045 0.085 5.295 1.105 ;
      RECT 5.905 0.085 6.235 1.105 ;
      RECT 6.835 0.085 7.165 1.105 ;
      RECT 7.765 0.085 8.095 1.105 ;
      RECT 8.695 0.085 9.025 1.105 ;
      RECT 9.625 0.085 9.955 1.105 ;
      RECT 10.555 0.085 10.885 1.105 ;
      RECT 11.555 0.085 11.885 1.13 ;
      RECT 10.14 2.02 10.47 2.98 ;
      RECT 10.125 1.92 10.47 2.02 ;
      RECT 10.125 0.35 10.375 1.92 ;
      RECT 9.19 2.02 9.52 2.98 ;
      RECT 9.195 1.92 9.52 2.02 ;
      RECT 9.195 0.35 9.445 1.92 ;
      RECT 8.24 2.02 8.57 2.98 ;
      RECT 8.265 1.92 8.57 2.02 ;
      RECT 8.265 0.35 8.515 1.92 ;
      RECT 7.34 1.92 7.67 2.98 ;
      RECT 7.34 0.35 7.585 1.92 ;
      RECT 6.44 2.02 6.77 2.98 ;
      RECT 6.42 1.92 6.77 2.02 ;
      RECT 6.42 0.35 6.655 1.92 ;
      RECT 5.54 2.02 5.87 2.98 ;
      RECT 5.51 1.92 5.87 2.02 ;
      RECT 5.51 0.35 5.725 1.92 ;
      RECT 4.64 2.02 4.97 2.98 ;
      RECT 4.615 1.92 4.97 2.02 ;
      RECT 4.615 0.35 4.865 1.92 ;
  END
END scs8ls_bufinv_16

MACRO scs8ls_bufinv_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 0.55 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.06 0.35 1.39 0.88 ;
        RECT 1.06 0.88 3.25 0.96 ;
        RECT 1.06 0.96 4.25 1.13 ;
        RECT 2.06 0.35 2.25 0.88 ;
        RECT 2.92 0.35 3.25 0.88 ;
        RECT 1.06 1.13 1.39 1.8 ;
        RECT 3.92 0.35 4.25 0.96 ;
        RECT 1.06 1.8 4.225 2.07 ;
    END
    ANTENNADIFFAREA 2.385 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 6.24 3.415 ;
      RECT 0.615 2.58 0.945 3.245 ;
      RECT 1.515 2.58 1.845 3.245 ;
      RECT 2.415 2.58 2.745 3.245 ;
      RECT 3.315 2.58 3.645 3.245 ;
      RECT 4.345 2.58 4.675 3.245 ;
      RECT 5.345 2.48 5.675 3.245 ;
      RECT 4.845 2.31 5.175 2.98 ;
      RECT 4.845 2.14 6.125 2.31 ;
      RECT 5.845 2.31 6.125 2.98 ;
      RECT 5.795 1.13 6.125 2.14 ;
      RECT 4.65 0.88 6.125 1.13 ;
      RECT 4.65 1.13 4.82 1.3 ;
      RECT 4.92 0.35 5.125 0.88 ;
      RECT 5.795 0.35 6.125 0.88 ;
      RECT 1.665 1.3 4.82 1.63 ;
      RECT 0 -0.085 6.24 0.085 ;
      RECT 4.42 0.085 4.75 0.71 ;
      RECT 5.295 0.085 5.625 0.71 ;
      RECT 0.56 0.085 0.89 0.84 ;
      RECT 1.56 0.085 1.89 0.71 ;
      RECT 2.42 0.085 2.75 0.71 ;
      RECT 3.42 0.085 3.75 0.79 ;
      RECT 0.115 2.24 4.565 2.41 ;
      RECT 4.395 1.97 4.565 2.24 ;
      RECT 4.395 1.8 5.605 1.97 ;
      RECT 4.99 1.32 5.605 1.8 ;
      RECT 0.115 2.41 0.445 2.98 ;
      RECT 0.115 1.95 0.445 2.24 ;
      RECT 0.72 1.18 0.89 2.24 ;
      RECT 0.13 1.01 0.89 1.18 ;
      RECT 0.13 0.35 0.38 1.01 ;
    LAYER mcon ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_bufinv_8

MACRO scs8ls_clkbuf_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475 0.35 1.805 0.79 ;
        RECT 1.565 0.79 1.805 1.82 ;
        RECT 1.345 1.82 1.805 2.98 ;
    END
    ANTENNADIFFAREA 0.4494 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.3 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.231 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.005 1.13 1.395 1.63 ;
      RECT 0.115 0.96 1.395 1.13 ;
      RECT 0.345 2.12 0.675 2.98 ;
      RECT 0.345 1.95 1.175 2.12 ;
      RECT 1.005 1.63 1.175 1.95 ;
      RECT 0.115 0.35 0.445 0.96 ;
      RECT 0 -0.085 1.92 0.085 ;
      RECT 0.615 0.085 1.305 0.68 ;
      RECT 0 3.245 1.92 3.415 ;
      RECT 0.845 2.29 1.175 3.245 ;
    LAYER mcon ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_clkbuf_1

MACRO scs8ls_clkbuf_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.795 1.78 ;
    END
    ANTENNAGATEAREA 0.924 ;
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2.39 1.92 9.09 2.15 ;
    END
    ANTENNADIFFAREA 3.6288 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 1.94 1.18 8.64 1.41 ;
    LAYER li1 ;
      RECT 8.225 1.19 8.555 1.52 ;
      RECT 7.295 1.19 7.625 1.52 ;
      RECT 6.365 1.19 6.695 1.52 ;
      RECT 5.425 1.19 5.755 1.52 ;
      RECT 4.51 1.19 4.84 1.52 ;
      RECT 3.67 1.19 4 1.52 ;
      RECT 2.835 1.19 3.105 1.52 ;
      RECT 7.84 1.86 8.05 2.98 ;
      RECT 7.795 1.69 8.05 1.86 ;
      RECT 7.795 0.35 8.045 1.69 ;
      RECT 0.115 0.085 0.365 0.81 ;
      RECT 0 -0.085 9.6 0.085 ;
      RECT 0.975 0.085 1.225 0.81 ;
      RECT 1.855 0.085 2.185 0.81 ;
      RECT 2.865 0.085 3.035 0.68 ;
      RECT 3.67 0.085 3.895 0.725 ;
      RECT 4.51 0.085 4.835 0.74 ;
      RECT 5.435 0.085 5.765 0.68 ;
      RECT 6.365 0.085 6.695 0.68 ;
      RECT 7.295 0.085 7.625 0.68 ;
      RECT 8.225 0.085 8.555 0.68 ;
      RECT 9.155 0.085 9.485 0.745 ;
      RECT 8.75 1.86 8.97 2.98 ;
      RECT 8.725 1.83 8.97 1.86 ;
      RECT 8.725 0.35 8.975 1.83 ;
      RECT 0 3.245 9.6 3.415 ;
      RECT 1.1 2.29 1.27 3.245 ;
      RECT 2 2.29 2.25 3.245 ;
      RECT 2.83 2.03 3.16 3.245 ;
      RECT 3.73 2.03 4.06 3.245 ;
      RECT 4.63 2.03 4.96 3.245 ;
      RECT 5.53 2.03 5.86 3.245 ;
      RECT 6.43 2.03 6.76 3.245 ;
      RECT 7.33 2.03 7.66 3.245 ;
      RECT 8.23 2.03 8.56 3.245 ;
      RECT 9.15 2.03 9.48 3.245 ;
      RECT 0.12 1.95 0.37 3.245 ;
      RECT 2.43 2.12 2.66 2.98 ;
      RECT 2.39 0.35 2.66 2.12 ;
      RECT 0.57 2.12 0.9 2.98 ;
      RECT 0.57 1.95 2.135 2.12 ;
      RECT 1.47 2.12 1.8 2.98 ;
      RECT 1.965 1.41 2.135 1.95 ;
      RECT 1.965 1.18 2.21 1.41 ;
      RECT 1.965 1.15 2.135 1.18 ;
      RECT 0.545 0.98 2.135 1.15 ;
      RECT 0.545 0.35 0.795 0.98 ;
      RECT 1.425 0.35 1.675 0.98 ;
      RECT 6.945 1.86 7.15 2.98 ;
      RECT 6.865 1.69 7.15 1.86 ;
      RECT 6.865 0.35 7.115 1.69 ;
      RECT 6.04 1.86 6.245 2.98 ;
      RECT 5.935 1.69 6.245 1.86 ;
      RECT 5.935 0.35 6.185 1.69 ;
      RECT 5.14 1.86 5.35 2.98 ;
      RECT 5.025 1.69 5.35 1.86 ;
      RECT 5.025 0.35 5.255 1.69 ;
      RECT 4.23 1.86 4.43 2.98 ;
      RECT 4.17 1.69 4.43 1.86 ;
      RECT 4.17 0.745 4.34 1.69 ;
      RECT 4.075 0.35 4.34 0.745 ;
      RECT 3.34 1.86 3.545 2.98 ;
      RECT 3.275 1.69 3.545 1.86 ;
      RECT 3.275 0.35 3.5 1.69 ;
    LAYER mcon ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.375 1.21 7.545 1.38 ;
      RECT 3.75 1.21 3.92 1.38 ;
      RECT 6.445 1.21 6.615 1.38 ;
      RECT 5.505 1.21 5.675 1.38 ;
      RECT 4.59 1.21 4.76 1.38 ;
      RECT 8.78 1.95 8.95 2.12 ;
      RECT 2.46 1.95 2.63 2.12 ;
      RECT 3.36 1.95 3.53 2.12 ;
      RECT 4.245 1.95 4.415 2.12 ;
      RECT 5.16 1.95 5.33 2.12 ;
      RECT 6.06 1.95 6.23 2.12 ;
      RECT 6.96 1.95 7.13 2.12 ;
      RECT 7.86 1.95 8.03 2.12 ;
      RECT 8.305 1.21 8.475 1.38 ;
      RECT 2.01 1.21 2.18 1.38 ;
      RECT 2.89 1.21 3.06 1.38 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
  END
END scs8ls_clkbuf_16

MACRO scs8ls_clkbuf_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.01 1.495 2.15 ;
    END
    ANTENNAGATEAREA 0.231 ;
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 0.35 0.885 0.79 ;
        RECT 0.715 0.79 0.885 1.82 ;
        RECT 0.555 1.82 0.885 2.15 ;
    END
    ANTENNADIFFAREA 0.4536 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.535 2.49 1.835 2.98 ;
      RECT 0.215 2.32 1.835 2.49 ;
      RECT 1.665 0.81 1.835 2.32 ;
      RECT 1.475 0.35 1.835 0.81 ;
      RECT 0.215 1.63 0.385 2.32 ;
      RECT 0.215 0.96 0.545 1.63 ;
      RECT 0 3.245 1.92 3.415 ;
      RECT 0.105 2.66 0.435 3.245 ;
      RECT 1.005 2.66 1.335 3.245 ;
      RECT 0 -0.085 1.92 0.085 ;
      RECT 1.055 0.085 1.305 0.81 ;
      RECT 0.115 0.085 0.365 0.79 ;
    LAYER mcon ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_clkbuf_2

MACRO scs8ls_clkbuf_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.56 0.35 0.89 0.98 ;
        RECT 0.535 0.98 1.75 1.15 ;
        RECT 0.535 1.15 0.705 1.92 ;
        RECT 1.42 0.35 1.75 0.98 ;
        RECT 0.535 1.92 1.795 2.09 ;
        RECT 0.535 2.09 0.815 2.98 ;
        RECT 1.465 2.09 1.795 2.98 ;
    END
    ANTENNADIFFAREA 0.924 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.055 1.08 2.455 1.41 ;
    END
    ANTENNAGATEAREA 0.231 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.415 1.75 2.795 2.98 ;
      RECT 0.875 1.58 2.795 1.75 ;
      RECT 2.625 0.81 2.795 1.58 ;
      RECT 2.42 0.48 2.795 0.81 ;
      RECT 0.875 1.35 1.885 1.58 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 1.995 1.92 2.245 3.245 ;
      RECT 0.115 1.82 0.365 3.245 ;
      RECT 1.015 2.26 1.265 3.245 ;
      RECT 0 -0.085 2.88 0.085 ;
      RECT 1.92 0.085 2.25 0.81 ;
      RECT 0.13 0.085 0.38 0.81 ;
      RECT 1.07 0.085 1.24 0.81 ;
    LAYER mcon ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_clkbuf_4

MACRO scs8ls_a31o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.255 2.815 0.64 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.49 2.405 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535 1.49 1.865 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995 1.49 1.325 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A3

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.85 0.435 2.98 ;
        RECT 0.085 1.18 0.255 1.85 ;
        RECT 0.085 0.48 0.45 1.18 ;
    END
    ANTENNADIFFAREA 0.5041 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.79 0.81 3.155 0.98 ;
      RECT 2.985 0.085 3.155 0.81 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 0.62 0.085 1.2 0.98 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 1.735 2.31 2.145 3.245 ;
      RECT 0.605 1.97 1.065 3.245 ;
      RECT 0.62 1.15 3.095 1.32 ;
      RECT 2.845 1.32 3.095 2.98 ;
      RECT 2.28 0.81 2.61 1.15 ;
      RECT 0.425 1.35 0.825 1.68 ;
      RECT 0.62 1.32 0.825 1.35 ;
      RECT 1.235 2.14 1.565 2.98 ;
      RECT 1.235 1.97 2.645 2.14 ;
      RECT 2.315 2.14 2.645 2.98 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a31o_1

MACRO scs8ls_a31o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.82 0.92 2.98 ;
        RECT 0.615 1.13 0.785 1.82 ;
        RECT 0.615 0.35 0.89 1.13 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.18 3.735 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.18 1.855 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.18 2.425 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.665 1.18 3.235 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.385 1.89 3.725 2.86 ;
      RECT 1.135 1.72 3.725 1.89 ;
      RECT 1.135 0.84 3.18 1.01 ;
      RECT 2.85 0.35 3.18 0.84 ;
      RECT 1.135 1.63 1.305 1.72 ;
      RECT 0.955 1.3 1.305 1.63 ;
      RECT 1.135 1.01 1.305 1.3 ;
      RECT 1.795 2.23 2.125 2.86 ;
      RECT 1.795 2.06 3.215 2.23 ;
      RECT 2.885 2.23 3.215 2.86 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 2.35 2.4 2.68 3.245 ;
      RECT 1.09 2.06 1.625 3.245 ;
      RECT 0.185 1.82 0.435 3.245 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 1.06 0.085 1.73 0.6 ;
      RECT 3.36 0.085 3.69 1.01 ;
      RECT 0.115 0.085 0.445 1.13 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_a31o_2

MACRO scs8ls_a31o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.55 0.895 1.72 ;
        RECT 0.565 1.72 1.895 1.89 ;
        RECT 0.615 1 0.865 1.55 ;
        RECT 0.565 1.89 0.895 2.98 ;
        RECT 1.565 1.89 1.895 2.98 ;
        RECT 0.615 0.83 1.725 1 ;
        RECT 0.615 0.35 0.865 0.83 ;
        RECT 1.555 0.33 1.725 0.83 ;
    END
    ANTENNADIFFAREA 1.1382 ;
  END X

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.565 1.47 3.235 1.8 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.115 1.45 7.075 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.45 5.865 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.45 4.675 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 4.98 1.11 7.03 1.28 ;
      RECT 4.98 0.595 5.23 1.11 ;
      RECT 5.92 0.35 6.09 1.11 ;
      RECT 6.78 0.35 7.03 1.11 ;
      RECT 1.065 1.22 4.75 1.28 ;
      RECT 1.895 1.13 4.75 1.22 ;
      RECT 3.42 1.11 4.75 1.13 ;
      RECT 4.42 0.595 4.75 1.11 ;
      RECT 3.125 1.97 3.575 2.64 ;
      RECT 3.405 1.3 3.575 1.97 ;
      RECT 1.065 1.28 3.59 1.3 ;
      RECT 2.49 0.35 2.74 1.13 ;
      RECT 3.42 0.35 3.75 1.11 ;
      RECT 1.065 1.3 2.335 1.55 ;
      RECT 3.92 0.425 4.25 0.94 ;
      RECT 3.92 0.255 5.74 0.425 ;
      RECT 5.41 0.425 5.74 0.94 ;
      RECT 2.625 2.81 4.075 2.98 ;
      RECT 3.745 2.12 4.075 2.81 ;
      RECT 2.625 1.97 2.955 2.81 ;
      RECT 3.745 1.95 7.085 2.12 ;
      RECT 4.745 2.12 5.075 2.98 ;
      RECT 5.755 2.12 6.085 2.98 ;
      RECT 6.755 2.12 7.085 2.98 ;
      RECT 0 3.245 7.2 3.415 ;
      RECT 4.245 2.29 4.575 3.245 ;
      RECT 5.245 2.29 5.575 3.245 ;
      RECT 6.255 2.29 6.585 3.245 ;
      RECT 2.065 1.82 2.395 3.245 ;
      RECT 0.115 1.82 0.365 3.245 ;
      RECT 1.065 2.06 1.395 3.245 ;
      RECT 0 -0.085 7.2 0.085 ;
      RECT 1.93 0.085 2.26 0.96 ;
      RECT 2.92 0.085 3.25 0.96 ;
      RECT 6.27 0.085 6.6 0.94 ;
      RECT 0.115 0.085 0.445 1.13 ;
      RECT 1.045 0.085 1.375 0.66 ;
    LAYER mcon ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
  END
END scs8ls_a31o_4

MACRO scs8ls_a31oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535 1.18 1.865 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 0.81 1.315 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.18 2.775 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.455 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A3

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.255 1.89 2.755 2.98 ;
        RECT 0.625 1.72 2.755 1.89 ;
        RECT 0.625 0.52 0.795 1.72 ;
        RECT 0.625 0.35 2.06 0.52 ;
        RECT 1.73 0.52 2.06 1.01 ;
    END
    ANTENNADIFFAREA 0.6412 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.665 2.23 0.995 2.98 ;
      RECT 0.665 2.06 2.085 2.23 ;
      RECT 1.755 2.23 2.085 2.98 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 0.125 1.82 0.455 3.245 ;
      RECT 1.205 2.4 1.535 3.245 ;
      RECT 0 -0.085 2.88 0.085 ;
      RECT 2.23 0.085 2.56 1.01 ;
      RECT 0.125 0.085 0.455 1.01 ;
    LAYER mcon ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_a31oi_1

MACRO scs8ls_a31oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325 1.18 2.995 1.55 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.875 0.425 4.205 1.09 ;
        RECT 3.165 1.09 4.205 1.26 ;
        RECT 2.545 0.255 4.205 0.425 ;
        RECT 3.165 1.26 3.335 1.72 ;
        RECT 2.545 0.425 3.26 0.58 ;
        RECT 2.475 1.72 3.335 1.89 ;
        RECT 2.475 1.89 2.805 2.735 ;
    END
    ANTENNADIFFAREA 1.0908 ;
  END Y

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.26 0.435 1.55 ;
        RECT 0.105 1.09 2.115 1.26 ;
        RECT 1.785 1.26 2.115 1.55 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A3

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.505 1.43 4.195 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.43 1.545 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.045 0.75 3.705 0.92 ;
      RECT 3.43 0.67 3.705 0.75 ;
      RECT 1.045 0.595 1.375 0.75 ;
      RECT 0.545 0.425 0.875 0.92 ;
      RECT 0.545 0.255 1.875 0.425 ;
      RECT 1.545 0.425 1.875 0.58 ;
      RECT 2.015 2.905 3.255 3.075 ;
      RECT 2.975 2.23 3.255 2.905 ;
      RECT 2.975 2.06 4.205 2.23 ;
      RECT 3.925 2.23 4.205 2.98 ;
      RECT 3.875 1.95 4.205 2.06 ;
      RECT 2.015 2.12 2.275 2.905 ;
      RECT 0.115 1.95 2.275 2.12 ;
      RECT 0.115 2.12 0.365 2.98 ;
      RECT 1.065 2.12 1.395 2.98 ;
      RECT 0.115 1.82 0.365 1.95 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 3.425 2.4 3.755 3.245 ;
      RECT 0.565 2.29 0.895 3.245 ;
      RECT 1.595 2.29 1.845 3.245 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 0.115 0.085 0.365 0.92 ;
      RECT 2.045 0.085 2.375 0.58 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_a31oi_2

MACRO scs8ls_a31oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.18 4.69 1.95 ;
        RECT 4.445 1.95 8.075 2.12 ;
        RECT 4.445 1.13 8.525 1.18 ;
        RECT 6.845 2.12 7.175 2.735 ;
        RECT 7.745 2.12 8.075 2.735 ;
        RECT 4.35 1.01 8.525 1.13 ;
        RECT 4.35 0.965 5.84 1.01 ;
        RECT 6.51 0.35 6.84 1.01 ;
        RECT 8.195 0.35 8.525 1.01 ;
        RECT 4.35 0.77 4.685 0.965 ;
        RECT 5.51 0.595 5.84 0.965 ;
    END
    ANTENNADIFFAREA 1.62135 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.35 6.115 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415 1.35 4.195 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.745 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.35 8.515 1.78 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END B1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 6.345 2.905 8.525 3.075 ;
      RECT 8.255 1.95 8.525 2.905 ;
      RECT 3.865 2.46 4.195 2.98 ;
      RECT 3.865 2.12 4.195 2.29 ;
      RECT 0.115 1.95 4.195 2.12 ;
      RECT 0.115 2.12 0.395 2.98 ;
      RECT 1.065 2.12 1.295 2.935 ;
      RECT 1.965 2.12 3.195 2.15 ;
      RECT 1.915 1.82 2.245 1.95 ;
      RECT 1.965 2.15 2.195 2.95 ;
      RECT 2.865 2.15 3.195 2.98 ;
      RECT 3.865 2.29 6.675 2.46 ;
      RECT 4.865 2.46 5.675 2.93 ;
      RECT 6.345 2.46 6.675 2.905 ;
      RECT 7.375 2.29 7.575 2.905 ;
      RECT 2.35 0.255 6.34 0.425 ;
      RECT 6.01 0.425 6.34 0.84 ;
      RECT 2.35 0.425 2.655 0.84 ;
      RECT 3.29 0.425 3.62 0.84 ;
      RECT 4.935 0.425 5.265 0.795 ;
      RECT 0.13 1.01 4.12 1.18 ;
      RECT 2.825 0.595 3.12 1.01 ;
      RECT 3.79 0.595 4.12 1.01 ;
      RECT 0.13 0.35 0.38 1.01 ;
      RECT 1.07 0.35 1.24 1.01 ;
      RECT 1.92 0.33 2.17 1.01 ;
      RECT 0 -0.085 8.64 0.085 ;
      RECT 0.56 0.085 0.89 0.84 ;
      RECT 1.42 0.085 1.75 0.84 ;
      RECT 7.01 0.085 8.025 0.84 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 4.365 2.63 4.695 3.245 ;
      RECT 5.845 2.63 6.175 3.245 ;
      RECT 2.365 2.32 2.695 3.245 ;
      RECT 0.565 2.29 0.895 3.245 ;
      RECT 1.465 2.29 1.795 3.245 ;
      RECT 3.365 2.29 3.695 3.245 ;
    LAYER mcon ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
  END
END scs8ls_a31oi_4

MACRO scs8ls_a32o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.19 1.315 1.55 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A3

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.19 2.375 1.55 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.19 1.835 1.55 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.545 1.19 3.005 1.55 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.29 1.21 3.715 1.55 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B2

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.35 0.445 1.13 ;
        RECT 0.085 1.13 0.255 1.82 ;
        RECT 0.085 1.82 0.455 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.395 2.905 3.725 3.075 ;
      RECT 2.395 2.23 2.725 2.905 ;
      RECT 3.395 1.82 3.725 2.905 ;
      RECT 1.205 2.06 2.725 2.23 ;
      RECT 1.205 2.23 1.535 2.86 ;
      RECT 2.895 1.89 3.225 2.735 ;
      RECT 0.625 1.72 3.225 1.89 ;
      RECT 0.625 0.85 2.88 1.02 ;
      RECT 2.2 0.43 2.88 0.85 ;
      RECT 0.625 1.63 0.795 1.72 ;
      RECT 0.425 1.3 0.795 1.63 ;
      RECT 0.625 1.02 0.795 1.3 ;
      RECT 0.65 0.085 1.05 0.68 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 3.37 0.085 3.7 1.04 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 1.8 2.4 2.13 3.245 ;
      RECT 0.625 2.06 1.015 3.245 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a32o_1

MACRO scs8ls_a32o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.82 0.935 2.15 ;
        RECT 0.725 1.15 0.935 1.82 ;
        RECT 0.615 0.33 0.935 1.15 ;
    END
    ANTENNADIFFAREA 0.5506 ;
  END X

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.35 2.915 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.015 1.35 2.345 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445 1.35 1.775 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.155 1.35 3.715 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885 1.3 4.215 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.105 1.95 3.705 2.12 ;
      RECT 3.375 2.12 3.705 2.735 ;
      RECT 1.105 1.01 3.105 1.18 ;
      RECT 2.775 0.35 3.105 1.01 ;
      RECT 0.225 2.32 1.275 2.49 ;
      RECT 1.105 2.12 1.275 2.32 ;
      RECT 1.105 1.18 1.275 1.95 ;
      RECT 0.225 1.65 0.395 2.32 ;
      RECT 0.225 1.32 0.555 1.65 ;
      RECT 2.875 2.905 4.205 3.075 ;
      RECT 2.875 2.46 3.205 2.905 ;
      RECT 3.875 1.95 4.205 2.905 ;
      RECT 1.715 2.29 3.205 2.46 ;
      RECT 1.715 2.46 2.045 2.86 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 1.185 0.085 1.515 0.84 ;
      RECT 3.85 0.085 4.18 1.13 ;
      RECT 0.115 0.085 0.445 1.13 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 0.115 2.66 0.445 3.245 ;
      RECT 1.1 2.66 1.51 3.245 ;
      RECT 2.265 2.63 2.645 3.245 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a32o_2

MACRO scs8ls_a32o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.44 1.47 5.35 1.79 ;
        RECT 5.18 1.79 5.35 1.95 ;
        RECT 5.18 1.95 6.595 2.12 ;
        RECT 6.425 1.77 6.595 1.95 ;
        RECT 6.425 1.44 6.825 1.77 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505 1.45 2.835 1.78 ;
        RECT 2.57 0.425 2.74 1.45 ;
        RECT 2.57 0.255 4.415 0.425 ;
        RECT 4.085 0.425 4.415 0.585 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B2

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.355 1.48 ;
        RECT 0.125 1.48 0.815 1.65 ;
        RECT 0.125 0.93 1.9 1.18 ;
        RECT 0.565 1.65 0.815 1.85 ;
        RECT 1.57 0.43 1.9 0.93 ;
        RECT 0.615 0.41 0.82 0.93 ;
        RECT 0.565 1.85 1.795 2.02 ;
        RECT 0.565 2.02 0.815 2.98 ;
        RECT 1.515 2.02 1.795 3 ;
    END
    ANTENNADIFFAREA 1.0975 ;
  END X

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.635 1.45 6.115 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.065 1.45 8.035 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.45 3.715 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 5.37 0.765 5.62 0.94 ;
      RECT 5.37 0.595 6.56 0.765 ;
      RECT 6.31 0.765 6.56 1.27 ;
      RECT 6.74 1.1 8.045 1.27 ;
      RECT 7.715 0.59 8.045 1.1 ;
      RECT 6.74 0.425 6.99 1.1 ;
      RECT 4.94 0.255 6.99 0.425 ;
      RECT 4.94 0.425 5.19 0.94 ;
      RECT 2.91 0.925 3.24 1.21 ;
      RECT 2.91 0.755 4.18 0.925 ;
      RECT 2.91 0.595 3.24 0.755 ;
      RECT 4.595 2.29 7.095 2.46 ;
      RECT 5.785 2.46 6.115 2.9 ;
      RECT 6.815 2.46 7.095 3 ;
      RECT 6.765 2.12 7.095 2.29 ;
      RECT 6.765 1.95 8.045 2.12 ;
      RECT 7.715 2.12 8.045 2.98 ;
      RECT 2.525 2.905 4.925 3.075 ;
      RECT 4.595 2.46 4.925 2.905 ;
      RECT 2.525 2.29 2.855 2.905 ;
      RECT 3.525 2.29 3.855 2.905 ;
      RECT 4.595 1.96 4.925 2.29 ;
      RECT 3.42 1.11 6.13 1.28 ;
      RECT 5.8 0.935 6.13 1.11 ;
      RECT 3.025 2.12 3.355 2.735 ;
      RECT 2.015 1.95 4.355 2.12 ;
      RECT 4.025 2.12 4.355 2.735 ;
      RECT 3.885 1.28 4.055 1.95 ;
      RECT 3.42 1.095 3.75 1.11 ;
      RECT 2.015 1.68 2.185 1.95 ;
      RECT 0.985 1.35 2.185 1.68 ;
      RECT 4.35 0.755 4.755 0.94 ;
      RECT 4.585 0.085 4.755 0.755 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 7.19 0.085 7.545 0.92 ;
      RECT 2.07 0.085 2.4 1.18 ;
      RECT 0.115 0.085 0.445 0.76 ;
      RECT 0.99 0.085 1.4 0.76 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 6.285 2.63 6.645 3.245 ;
      RECT 7.265 2.29 7.545 3.245 ;
      RECT 1.965 2.29 2.295 3.245 ;
      RECT 0.115 1.82 0.365 3.245 ;
      RECT 1.015 2.19 1.345 3.245 ;
      RECT 5.21 2.63 5.615 3.245 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
  END
END scs8ls_a32o_4

MACRO scs8ls_a32oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.18 1.855 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.59 1.89 2.275 2.15 ;
        RECT 0.615 1.72 2.275 1.89 ;
        RECT 0.615 1.89 0.945 2.735 ;
        RECT 0.615 1.01 0.785 1.72 ;
        RECT 0.615 0.35 1.83 1.01 ;
    END
    ANTENNADIFFAREA 0.9988 ;
  END Y

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 0.44 2.525 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955 1.18 1.315 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.18 0.445 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.765 1.18 3.235 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A3

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.115 2.32 2.795 2.49 ;
      RECT 2.515 2.49 2.795 2.98 ;
      RECT 2.465 1.82 2.795 2.32 ;
      RECT 0.115 1.82 0.445 2.905 ;
      RECT 0.115 2.905 1.445 3.075 ;
      RECT 1.115 2.49 1.445 2.905 ;
      RECT 1.115 2.06 1.42 2.32 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 1.675 2.66 2.345 3.245 ;
      RECT 2.995 1.82 3.245 3.245 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.89 0.085 3.22 1.01 ;
      RECT 0.115 0.085 0.445 1.01 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_a32oi_1

MACRO scs8ls_a32oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.235 3.235 1.72 ;
        RECT 1.615 1.72 3.235 1.8 ;
        RECT 3.005 1.01 3.205 1.235 ;
        RECT 0.615 1.8 3.235 1.89 ;
        RECT 1.455 0.84 3.205 1.01 ;
        RECT 0.615 1.89 1.945 1.97 ;
        RECT 1.455 0.595 1.785 0.84 ;
        RECT 3.015 0.595 3.205 0.84 ;
        RECT 0.615 1.97 0.945 2.735 ;
        RECT 1.615 1.97 1.945 2.735 ;
    END
    ANTENNADIFFAREA 1.1928 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.18 2.775 1.55 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.35 4.375 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.785 1.18 6.115 1.55 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.18 2.275 1.55 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.63 0.355 1.78 ;
        RECT 0.125 1.3 1.09 1.63 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 6.24 3.415 ;
      RECT 2.57 2.4 3.28 3.245 ;
      RECT 3.905 2.29 4.25 3.245 ;
      RECT 5.045 2.06 5.375 3.245 ;
      RECT 0 -0.085 6.24 0.085 ;
      RECT 4.935 0.085 5.185 0.84 ;
      RECT 5.795 0.085 6.125 1.01 ;
      RECT 0.545 0.085 0.875 0.79 ;
      RECT 2.115 2.12 3.735 2.23 ;
      RECT 3.45 2.23 3.735 2.98 ;
      RECT 2.115 2.06 4.875 2.12 ;
      RECT 4.42 2.12 4.875 2.98 ;
      RECT 3.405 1.95 4.875 2.06 ;
      RECT 4.545 1.89 4.875 1.95 ;
      RECT 4.545 1.72 5.875 1.89 ;
      RECT 5.545 1.89 5.875 2.98 ;
      RECT 0.115 2.905 2.4 3.075 ;
      RECT 2.115 2.23 2.4 2.905 ;
      RECT 0.115 1.95 0.445 2.905 ;
      RECT 1.115 2.14 1.445 2.905 ;
      RECT 2.515 0.255 4.705 0.425 ;
      RECT 3.375 0.425 3.705 1.13 ;
      RECT 4.375 0.425 4.705 0.84 ;
      RECT 2.515 0.425 2.845 0.67 ;
      RECT 3.875 1.01 5.615 1.18 ;
      RECT 3.875 0.595 4.205 1.01 ;
      RECT 5.365 0.35 5.615 1.01 ;
      RECT 1.105 0.255 2.285 0.425 ;
      RECT 1.955 0.425 2.285 0.67 ;
      RECT 0.115 0.96 1.275 1.13 ;
      RECT 1.105 0.425 1.275 0.96 ;
      RECT 0.115 0.35 0.365 0.96 ;
    LAYER mcon ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_a32oi_2

MACRO scs8ls_a32oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.82 0.77 6.35 1.01 ;
        RECT 2.4 1.01 6.35 1.13 ;
        RECT 6.18 1.13 6.35 1.95 ;
        RECT 2.4 1.13 5.15 1.18 ;
        RECT 2.4 0.88 3.66 1.01 ;
        RECT 0.615 1.95 6.35 2.12 ;
        RECT 2.4 0.595 2.73 0.88 ;
        RECT 0.615 2.12 0.945 2.735 ;
        RECT 1.515 2.12 1.845 2.735 ;
        RECT 2.515 2.12 2.845 2.735 ;
        RECT 3.515 2.12 3.845 2.735 ;
    END
    ANTENNADIFFAREA 2.387 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.35 5.805 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.735 1.35 8.515 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.765 1.35 10.435 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 4.195 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.795 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.115 2.905 4.345 3.075 ;
      RECT 4.015 2.46 4.345 2.905 ;
      RECT 4.015 2.29 7.435 2.46 ;
      RECT 5.105 2.46 5.435 2.98 ;
      RECT 6.105 2.46 6.435 2.98 ;
      RECT 7.105 2.46 7.435 2.98 ;
      RECT 7.105 2.12 7.435 2.29 ;
      RECT 7.105 1.95 10.44 2.12 ;
      RECT 8.105 2.12 8.435 2.98 ;
      RECT 9.105 2.12 9.435 2.98 ;
      RECT 10.11 2.12 10.44 2.98 ;
      RECT 0.115 1.95 0.445 2.905 ;
      RECT 1.145 2.29 1.315 2.905 ;
      RECT 2.015 2.29 2.345 2.905 ;
      RECT 3.015 2.29 3.345 2.905 ;
      RECT 6.54 1.01 9.935 1.18 ;
      RECT 6.54 0.85 7.735 1.01 ;
      RECT 8.905 0.35 9.075 1.01 ;
      RECT 9.765 0.35 9.935 1.01 ;
      RECT 6.54 0.77 6.87 0.85 ;
      RECT 4.32 0.35 8.165 0.6 ;
      RECT 7.835 0.6 8.165 0.68 ;
      RECT 4.32 0.6 4.65 0.84 ;
      RECT 2.05 0.255 4.09 0.425 ;
      RECT 2.9 0.425 3.23 0.71 ;
      RECT 3.76 0.425 4.09 0.71 ;
      RECT 0.115 1.01 2.22 1.18 ;
      RECT 2.05 0.425 2.22 1.01 ;
      RECT 0.115 0.35 0.445 1.01 ;
      RECT 1.125 0.35 1.295 1.01 ;
      RECT 0 3.245 10.56 3.415 ;
      RECT 4.605 2.63 4.935 3.245 ;
      RECT 5.605 2.63 5.935 3.245 ;
      RECT 6.605 2.63 6.935 3.245 ;
      RECT 7.605 2.29 7.935 3.245 ;
      RECT 8.605 2.29 8.935 3.245 ;
      RECT 9.605 2.29 9.935 3.245 ;
      RECT 0 -0.085 10.56 0.085 ;
      RECT 8.395 0.085 8.725 0.84 ;
      RECT 9.255 0.085 9.585 0.84 ;
      RECT 10.115 0.085 10.445 1.13 ;
      RECT 0.615 0.085 0.945 0.84 ;
      RECT 1.475 0.085 1.805 0.84 ;
    LAYER mcon ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
  END
END scs8ls_a32oi_4

MACRO scs8ls_a41o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.29 1.12 0.94 ;
        RECT 0.115 0.94 0.355 1.82 ;
        RECT 0.115 1.82 0.445 2.98 ;
    END
    ANTENNADIFFAREA 1.0408 ;
  END X

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.45 1.815 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.135 1.18 3.715 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 0.44 2.895 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025 1.45 2.355 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885 1.18 4.215 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A4

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.575 1.11 2.12 1.28 ;
      RECT 1.79 0.35 2.12 1.11 ;
      RECT 1.145 1.95 1.635 2.98 ;
      RECT 1.145 1.55 1.315 1.95 ;
      RECT 0.575 1.28 1.315 1.55 ;
      RECT 1.805 2.12 2.135 2.98 ;
      RECT 1.805 1.95 3.165 2.12 ;
      RECT 2.835 2.12 3.165 2.98 ;
      RECT 2.835 1.89 3.165 1.95 ;
      RECT 2.835 1.72 4.185 1.89 ;
      RECT 3.855 1.89 4.185 2.98 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 2.305 2.29 2.635 3.245 ;
      RECT 3.335 2.06 3.665 3.245 ;
      RECT 0.645 1.82 0.895 3.245 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 3.83 0.085 4.16 1.01 ;
      RECT 1.29 0.085 1.62 0.94 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_a41o_1

MACRO scs8ls_a41o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385 0.35 3.715 0.77 ;
        RECT 3.385 0.77 4.185 0.94 ;
        RECT 4.015 0.94 4.185 1.82 ;
        RECT 3.855 1.82 4.185 2.98 ;
    END
    ANTENNADIFFAREA 0.6394 ;
  END X

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.45 2.925 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.455 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.845 0.44 1.315 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 0.44 1.815 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025 1.45 2.355 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.095 1.28 3.845 1.55 ;
      RECT 2.23 1.11 3.845 1.28 ;
      RECT 2.795 2.12 3.125 2.98 ;
      RECT 2.795 1.95 3.265 2.12 ;
      RECT 3.095 1.55 3.265 1.95 ;
      RECT 2.23 0.35 2.56 1.11 ;
      RECT 1.115 1.95 2.625 2.12 ;
      RECT 2.295 2.12 2.625 2.98 ;
      RECT 1.115 2.12 1.445 2.98 ;
      RECT 1.115 1.89 1.445 1.95 ;
      RECT 0.115 1.72 1.445 1.89 ;
      RECT 0.115 1.89 0.445 2.98 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 4.355 1.82 4.685 3.245 ;
      RECT 1.615 2.29 2.125 3.245 ;
      RECT 3.355 2.27 3.685 3.245 ;
      RECT 0.615 2.06 0.945 3.245 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 3.885 0.085 4.685 0.6 ;
      RECT 2.79 0.085 3.12 0.94 ;
      RECT 0.15 0.085 0.48 1.01 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_a41o_2

MACRO scs8ls_a41o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.45 0.55 1.78 ;
    END
    ANTENNAGATEAREA 0.522 ;
  END B1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.9 1.45 5.635 1.78 ;
    END
    ANTENNAGATEAREA 0.522 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.45 4.195 1.78 ;
    END
    ANTENNAGATEAREA 0.522 ;
  END A1

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.325 1.45 8.035 1.78 ;
    END
    ANTENNAGATEAREA 0.522 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.45 7.075 1.78 ;
    END
    ANTENNAGATEAREA 0.522 ;
  END A3

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555 1.17 3.305 1.84 ;
        RECT 2.075 1.84 3.305 2.12 ;
        RECT 1.55 1 3.305 1.17 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 6.86 1.11 8.05 1.28 ;
      RECT 6.86 0.425 7.11 1.11 ;
      RECT 7.79 0.35 8.05 1.11 ;
      RECT 6 0.255 7.11 0.425 ;
      RECT 6 0.425 6.33 0.94 ;
      RECT 1.065 2.29 4.375 2.46 ;
      RECT 4.045 2.46 4.375 2.98 ;
      RECT 4.045 2.12 4.375 2.29 ;
      RECT 4.045 1.95 7.595 2.12 ;
      RECT 5.265 2.12 5.595 2.98 ;
      RECT 6.265 2.12 6.595 2.98 ;
      RECT 7.265 2.12 7.595 2.98 ;
      RECT 0.115 2.905 1.395 3.075 ;
      RECT 1.065 2.46 1.395 2.905 ;
      RECT 0.115 1.95 0.445 2.905 ;
      RECT 1.065 1.94 1.395 2.29 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 3.425 2.65 3.775 3.245 ;
      RECT 2.525 2.63 2.855 3.245 ;
      RECT 4.635 2.29 5.095 3.245 ;
      RECT 5.765 2.29 6.095 3.245 ;
      RECT 6.765 2.29 7.095 3.245 ;
      RECT 7.795 1.95 8.045 3.245 ;
      RECT 1.625 2.63 1.955 3.245 ;
      RECT 5.025 1.11 6.68 1.28 ;
      RECT 5.025 0.77 5.285 1.11 ;
      RECT 6.51 0.595 6.68 1.11 ;
      RECT 3.815 0.77 4.845 1.15 ;
      RECT 3.815 0.7 3.985 0.77 ;
      RECT 4.675 0.6 4.845 0.77 ;
      RECT 4.675 0.33 5.785 0.6 ;
      RECT 5.455 0.6 5.785 0.94 ;
      RECT 0.54 0.66 3.645 0.83 ;
      RECT 3.475 0.425 3.645 0.66 ;
      RECT 3.475 0.255 4.495 0.425 ;
      RECT 4.165 0.425 4.495 0.6 ;
      RECT 0.615 1.95 0.89 2.735 ;
      RECT 0.72 1.67 0.89 1.95 ;
      RECT 0.72 1.25 1.225 1.34 ;
      RECT 0.54 0.83 1.225 1.25 ;
      RECT 0.54 0.47 0.87 0.66 ;
      RECT 0.72 1.34 2.385 1.67 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 3.055 0.085 3.305 0.49 ;
      RECT 7.29 0.085 7.62 0.94 ;
      RECT 0.11 0.085 0.36 1.25 ;
      RECT 1.045 0.085 1.375 0.49 ;
      RECT 2.055 0.085 2.385 0.49 ;
    LAYER mcon ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a41o_4

MACRO scs8ls_a41oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.35 1.955 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.35 1.335 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A4

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.3 0.435 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.3 3.255 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.195 1.35 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.13 0.835 1.95 ;
        RECT 0.115 1.95 0.835 2.12 ;
        RECT 0.115 0.96 3.22 1.13 ;
        RECT 0.115 2.12 0.445 2.98 ;
        RECT 0.115 0.35 0.445 0.96 ;
        RECT 2.89 0.35 3.22 0.96 ;
    END
    ANTENNADIFFAREA 0.7522 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.615 2.46 0.945 2.98 ;
      RECT 0.615 2.29 1.275 2.46 ;
      RECT 1.105 1.95 3.245 2.29 ;
      RECT 2.915 2.29 3.245 2.98 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 1.115 2.63 1.785 3.245 ;
      RECT 2.405 2.46 2.745 3.245 ;
      RECT 1.445 2.46 1.785 2.63 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 0.615 0.085 1.26 0.68 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_a41oi_1

MACRO scs8ls_a41oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.085 1.78 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END B1

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.35 5.635 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.35 4.675 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.63 3.715 1.78 ;
        RECT 2.665 1.3 3.715 1.63 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965 1.26 2.275 1.65 ;
        RECT 1.965 1.65 2.135 1.95 ;
        RECT 1.685 1.18 2.275 1.26 ;
        RECT 0.615 1.95 2.135 2.12 ;
        RECT 0.615 1.09 2.275 1.18 ;
        RECT 0.615 2.12 0.945 2.735 ;
        RECT 0.615 1.01 1.935 1.09 ;
        RECT 1.685 0.595 1.935 1.01 ;
        RECT 0.615 0.4 0.945 1.01 ;
    END
    ANTENNADIFFAREA 0.8101 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415 1.43 1.795 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 1.615 2.65 2.135 3.245 ;
      RECT 2.805 2.29 3.135 3.245 ;
      RECT 3.805 2.29 4.135 3.245 ;
      RECT 4.84 2.29 5.17 3.245 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 4.815 0.085 5.145 0.84 ;
      RECT 0.115 0.085 0.445 1.18 ;
      RECT 4.305 2.12 4.67 3 ;
      RECT 2.305 1.95 5.645 2.12 ;
      RECT 2.305 2.12 2.635 2.29 ;
      RECT 3.305 2.12 3.635 2.98 ;
      RECT 2.305 1.82 2.635 1.95 ;
      RECT 1.115 2.29 2.635 2.46 ;
      RECT 2.305 2.46 2.635 2.98 ;
      RECT 5.34 2.12 5.645 3 ;
      RECT 0.115 1.95 0.445 2.905 ;
      RECT 1.115 2.46 1.445 2.905 ;
      RECT 0.115 2.905 1.445 3.075 ;
      RECT 2.965 0.92 3.295 1.08 ;
      RECT 2.105 0.75 3.295 0.92 ;
      RECT 2.105 0.425 2.355 0.75 ;
      RECT 1.175 0.255 2.355 0.425 ;
      RECT 1.175 0.425 1.505 0.84 ;
      RECT 3.955 0.58 4.285 0.68 ;
      RECT 2.535 0.33 4.285 0.58 ;
      RECT 4.465 1.13 5.645 1.18 ;
      RECT 3.525 1.01 5.645 1.13 ;
      RECT 3.525 0.85 4.635 1.01 ;
      RECT 5.315 0.35 5.645 1.01 ;
      RECT 4.465 0.35 4.635 0.85 ;
    LAYER mcon ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_a41oi_2

MACRO scs8ls_a41oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.43 1.78 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END B1

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285 1.35 9.955 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A4

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.35 8.035 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A3

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.65 4.675 1.78 ;
        RECT 3.965 1.32 5.62 1.65 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.285 1.35 3.295 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.465 1.55 3.715 1.95 ;
        RECT 0.615 1.95 3.715 2.12 ;
        RECT 3.465 1 3.635 1.55 ;
        RECT 0.615 2.12 0.945 2.735 ;
        RECT 1.645 2.12 1.815 2.735 ;
        RECT 1.645 1.82 2.105 1.95 ;
        RECT 3.305 0.595 3.635 1 ;
        RECT 1.815 1.18 2.105 1.82 ;
        RECT 0.545 1.01 2.435 1.18 ;
        RECT 2.105 0.595 2.435 1.01 ;
        RECT 0.545 0.35 0.875 1.01 ;
    END
    ANTENNADIFFAREA 1.4476 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.805 0.62 4.135 1.13 ;
      RECT 3.805 0.425 5.925 0.62 ;
      RECT 1.605 0.255 5.925 0.425 ;
      RECT 1.605 0.425 1.935 0.84 ;
      RECT 2.605 0.425 3.135 1.13 ;
      RECT 4.305 0.79 7.775 1.13 ;
      RECT 7.445 0.77 7.775 0.79 ;
      RECT 7.955 1.01 9.965 1.18 ;
      RECT 7.955 0.6 8.125 1.01 ;
      RECT 8.815 0.35 8.985 1.01 ;
      RECT 9.715 0.35 9.965 1.01 ;
      RECT 6.155 0.35 8.125 0.6 ;
      RECT 6.155 0.6 6.485 0.62 ;
      RECT 2.015 2.29 4.3 2.46 ;
      RECT 3.97 2.46 4.3 2.98 ;
      RECT 3.97 2.12 4.3 2.29 ;
      RECT 3.97 1.95 9.96 2.12 ;
      RECT 4.93 2.12 5.26 2.98 ;
      RECT 5.88 2.12 6.21 2.98 ;
      RECT 6.83 2.12 7.16 2.98 ;
      RECT 7.78 2.12 8.11 2.98 ;
      RECT 8.73 2.12 9.06 2.98 ;
      RECT 9.63 2.12 9.96 2.98 ;
      RECT 4.93 1.82 5.26 1.95 ;
      RECT 0.115 1.95 0.445 2.905 ;
      RECT 1.115 2.29 1.445 2.905 ;
      RECT 0.115 2.905 2.345 3.075 ;
      RECT 2.015 2.46 2.345 2.905 ;
      RECT 3.015 2.46 3.345 2.98 ;
      RECT 0 3.245 10.08 3.415 ;
      RECT 2.515 2.63 2.845 3.245 ;
      RECT 3.545 2.63 3.795 3.245 ;
      RECT 4.5 2.29 4.75 3.245 ;
      RECT 5.46 2.29 5.71 3.245 ;
      RECT 6.41 2.29 6.66 3.245 ;
      RECT 7.36 2.29 7.61 3.245 ;
      RECT 8.28 2.29 8.53 3.245 ;
      RECT 9.26 2.29 9.43 3.245 ;
      RECT 0 -0.085 10.08 0.085 ;
      RECT 8.305 0.085 8.635 0.84 ;
      RECT 9.165 0.085 9.495 0.84 ;
      RECT 0.115 0.085 0.365 1.13 ;
      RECT 1.045 0.085 1.375 0.84 ;
    LAYER mcon ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
  END
END scs8ls_a41oi_4

MACRO scs8ls_and2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.92 1.85 2.315 2.98 ;
        RECT 2.145 1.18 2.315 1.85 ;
        RECT 1.84 0.47 2.315 1.18 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.075 1.18 1.405 1.68 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.255 0.835 0.67 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.58 1.35 1.975 1.68 ;
      RECT 0.855 2.02 1.185 3 ;
      RECT 0.26 1.85 1.75 2.02 ;
      RECT 1.58 1.68 1.75 1.85 ;
      RECT 0.26 0.84 0.59 1.85 ;
      RECT 0 3.245 2.4 3.415 ;
      RECT 0.35 2.19 0.685 3.245 ;
      RECT 1.39 2.19 1.72 3.245 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 1.34 0.085 1.67 1.01 ;
    LAYER mcon ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_and2_1

MACRO scs8ls_and2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.595 1.89 1.845 2.98 ;
        RECT 1.595 1.72 2.01 1.89 ;
        RECT 1.84 1.02 2.01 1.72 ;
        RECT 1.625 0.85 2.01 1.02 ;
        RECT 1.625 0.79 1.795 0.85 ;
        RECT 1.465 0.35 1.795 0.79 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.3 1.085 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.3 0.435 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.255 1.22 1.67 1.55 ;
      RECT 0.64 2.12 0.89 2.98 ;
      RECT 0.64 1.95 1.425 2.12 ;
      RECT 1.255 1.55 1.425 1.95 ;
      RECT 1.255 1.13 1.425 1.22 ;
      RECT 0.135 0.96 1.425 1.13 ;
      RECT 0.135 0.35 0.465 0.96 ;
      RECT 0 3.245 2.4 3.415 ;
      RECT 2.045 2.06 2.295 3.245 ;
      RECT 1.06 2.29 1.39 3.245 ;
      RECT 0.11 1.95 0.44 3.245 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 1.975 0.085 2.285 0.68 ;
      RECT 0.955 0.085 1.285 0.79 ;
    LAYER mcon ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_and2_2

MACRO scs8ls_and2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.255 1.345 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.444 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.45 3.255 1.78 ;
    END
    ANTENNAGATEAREA 0.444 ;
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.55 0.835 1.845 ;
        RECT 0.545 1.845 1.715 2.015 ;
        RECT 0.545 1.175 0.795 1.55 ;
        RECT 0.545 2.015 0.815 2.98 ;
        RECT 1.465 2.015 1.715 2.98 ;
        RECT 0.545 1.005 1.725 1.175 ;
        RECT 0.545 0.475 0.795 1.005 ;
        RECT 1.475 0.475 1.725 1.005 ;
    END
    ANTENNADIFFAREA 1.2198 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.495 0.425 2.825 1.175 ;
      RECT 2.495 0.255 3.675 0.425 ;
      RECT 3.505 0.425 3.675 0.94 ;
      RECT 1.885 1.95 3.67 2.12 ;
      RECT 3.5 2.12 3.67 2.905 ;
      RECT 3.5 1.28 3.67 1.95 ;
      RECT 2.995 1.11 3.67 1.28 ;
      RECT 2.995 0.595 3.325 1.11 ;
      RECT 2.47 2.12 2.8 2.905 ;
      RECT 1.885 1.675 2.055 1.95 ;
      RECT 1.005 1.345 2.055 1.675 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 1.935 2.29 2.265 3.245 ;
      RECT 2.97 2.29 3.3 3.245 ;
      RECT 3.87 2.025 4.2 3.245 ;
      RECT 0.115 1.82 0.365 3.245 ;
      RECT 1.015 2.185 1.265 3.245 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 1.985 0.085 2.315 1.175 ;
      RECT 3.875 0.085 4.205 1.255 ;
      RECT 0.115 0.085 0.365 1.255 ;
      RECT 0.975 0.085 1.305 0.835 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_and2_4

MACRO scs8ls_and2b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.77 1.82 3.255 2.98 ;
        RECT 3.085 1.15 3.255 1.82 ;
        RECT 2.915 0.37 3.255 1.15 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 0.55 2.15 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END AN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 2.375 1.78 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END B

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.115 2.32 1.165 2.65 ;
      RECT 0.81 1.18 1.14 2.32 ;
      RECT 0.115 1.01 1.14 1.18 ;
      RECT 0.115 0.35 0.445 1.01 ;
      RECT 2.575 1.32 2.915 1.65 ;
      RECT 1.705 1.95 2.065 2.7 ;
      RECT 1.31 0.98 2.745 1.15 ;
      RECT 2.575 1.15 2.745 1.32 ;
      RECT 1.705 1.15 1.875 1.95 ;
      RECT 1.31 0.47 1.64 0.98 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.27 1.95 2.6 3.245 ;
      RECT 1.365 1.82 1.535 3.245 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 0.615 0.085 0.945 0.84 ;
      RECT 2.13 0.085 2.745 0.81 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_and2b_1

MACRO scs8ls_and2b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 0.55 1.78 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END AN

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.18 2.525 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.82 1.515 2.15 ;
        RECT 1.115 1.13 1.285 1.82 ;
        RECT 1.115 0.35 1.445 1.13 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.685 1.87 2.795 2.15 ;
      RECT 1.685 0.84 3.22 1.01 ;
      RECT 2.89 1.01 3.22 1.13 ;
      RECT 2.89 0.35 3.22 0.84 ;
      RECT 1.685 1.63 1.855 1.87 ;
      RECT 1.455 1.3 1.855 1.63 ;
      RECT 1.685 1.01 1.855 1.3 ;
      RECT 0.115 2.32 3.135 2.49 ;
      RECT 2.965 1.63 3.135 2.32 ;
      RECT 2.765 1.3 3.135 1.63 ;
      RECT 0.115 2.49 0.445 2.7 ;
      RECT 0.115 1.95 0.89 2.32 ;
      RECT 0.72 1.18 0.89 1.95 ;
      RECT 0.115 1.01 0.89 1.18 ;
      RECT 0.115 0.35 0.445 1.01 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 0.65 2.66 0.98 3.245 ;
      RECT 1.635 2.66 2.26 3.245 ;
      RECT 2.915 2.66 3.245 3.245 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 1.615 0.085 2.4 0.6 ;
      RECT 0.615 0.085 0.945 0.84 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_and2b_2

MACRO scs8ls_and2b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.15 4.675 1.48 ;
        RECT 3.995 1.48 4.675 1.65 ;
        RECT 3.095 0.98 4.675 1.15 ;
        RECT 3.995 1.65 4.165 1.82 ;
        RECT 3.095 0.35 3.265 0.98 ;
        RECT 3.91 0.35 4.16 0.98 ;
        RECT 3.095 1.82 4.165 1.99 ;
        RECT 3.095 1.99 3.265 2.98 ;
        RECT 3.995 1.99 4.165 2.98 ;
    END
    ANTENNADIFFAREA 1.0938 ;
  END X

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.18 2.585 1.62 ;
        RECT 0.975 1.62 2.585 1.79 ;
        RECT 0.975 1.435 1.305 1.62 ;
    END
    ANTENNAGATEAREA 0.444 ;
  END B

  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.45 0.805 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END AN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.21 0.585 1.47 0.925 ;
      RECT 1.21 0.335 2.4 0.585 ;
      RECT 0.085 1.095 1.845 1.265 ;
      RECT 1.515 1.265 1.845 1.45 ;
      RECT 0.085 0.35 0.54 1.095 ;
      RECT 0.085 1.95 0.355 2.98 ;
      RECT 0.085 1.265 0.255 1.95 ;
      RECT 2.755 1.32 3.825 1.65 ;
      RECT 1.075 1.96 2.925 2.13 ;
      RECT 2.045 2.13 2.375 2.98 ;
      RECT 2.755 1.65 2.925 1.96 ;
      RECT 2.755 0.925 2.925 1.32 ;
      RECT 1.64 0.755 2.925 0.925 ;
      RECT 1.075 2.13 1.405 2.98 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 4.34 0.085 4.67 0.81 ;
      RECT 0.71 0.085 1.04 0.925 ;
      RECT 2.57 0.085 2.9 0.585 ;
      RECT 3.445 0.085 3.695 0.81 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 4.365 1.82 4.695 3.245 ;
      RECT 1.605 2.3 1.855 3.245 ;
      RECT 2.565 2.3 2.895 3.245 ;
      RECT 0.555 2.1 0.885 3.245 ;
      RECT 3.465 2.16 3.795 3.245 ;
    LAYER mcon ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_and2b_4

MACRO scs8ls_and3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.48 1.85 2.765 2.98 ;
        RECT 2.595 1.18 2.765 1.85 ;
        RECT 2.195 1.01 2.765 1.18 ;
        RECT 2.195 0.48 2.525 1.01 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.45 1.815 1.78 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END C

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.845 1.18 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.255 1.315 0.57 ;
        RECT 1.085 0.57 1.315 0.67 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.115 1.95 2.24 2.12 ;
      RECT 2.07 1.68 2.24 1.95 ;
      RECT 2.07 1.35 2.4 1.68 ;
      RECT 1.115 2.12 1.4 2.85 ;
      RECT 0.115 2.12 0.445 2.85 ;
      RECT 0.115 0.74 0.48 1.95 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 0.615 2.29 0.945 3.245 ;
      RECT 1.57 2.29 2.31 3.245 ;
      RECT 0 -0.085 2.88 0.085 ;
      RECT 1.695 0.085 2.025 1.18 ;
    LAYER mcon ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_and3_1

MACRO scs8ls_and3_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.905 1.18 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END B

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.255 1.315 0.67 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.18 0.81 2.755 1.17 ;
        RECT 2.555 1.17 2.725 1.84 ;
        RECT 2.18 0.39 2.51 0.81 ;
        RECT 2.375 1.84 2.725 2.98 ;
    END
    ANTENNADIFFAREA 0.5728 ;
  END X

  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.43 1.815 1.78 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END C

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.035 1.34 2.385 1.67 ;
      RECT 1.205 2.12 1.535 2.78 ;
      RECT 0.185 1.95 2.205 2.12 ;
      RECT 2.035 1.67 2.205 1.95 ;
      RECT 0.185 2.12 0.515 2.78 ;
      RECT 0.185 1.34 0.515 1.95 ;
      RECT 0.185 0.84 0.54 1.34 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.895 1.82 3.225 3.245 ;
      RECT 0.685 2.29 1.015 3.245 ;
      RECT 1.875 2.29 2.205 3.245 ;
      RECT 2.925 0.64 3.245 1.17 ;
      RECT 2.68 0.085 3.245 0.64 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 1.68 0.085 2.01 1.17 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_and3_2

MACRO scs8ls_a221o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435 0.255 1.765 0.565 ;
        RECT 1.595 0.565 1.765 1.04 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845 0.505 7.045 0.67 ;
        RECT 6.47 0.255 7.045 0.505 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B2

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 0.505 2.755 0.67 ;
        RECT 2.275 0.255 2.755 0.505 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.615 1.3 9.495 1.75 ;
        RECT 9.095 1.21 9.495 1.3 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405 1.47 5.735 2.15 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END C1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
    END
  END vpwr

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.095 1.225 3.265 1.365 ;
        RECT 2.975 1.365 3.265 1.41 ;
        RECT 2.975 1.18 3.265 1.225 ;
        RECT 0.095 1.365 0.385 1.41 ;
        RECT 0.095 1.18 0.385 1.225 ;
    END
    ANTENNADIFFAREA 1.0864 ;
    ANTENNAPARTIALMETALSIDEAREA 2.205 LAYER met1 ;
  END X

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.255 1.24 2.76 1.41 ;
      RECT 2.51 0.84 2.76 1.24 ;
      RECT 1.255 0.905 1.425 1.24 ;
      RECT 0.315 0.735 1.425 0.905 ;
      RECT 0.315 0.905 0.565 1.01 ;
      RECT 0.315 0.655 0.565 0.735 ;
      RECT 7.685 0.255 8.925 0.425 ;
      RECT 8.625 0.425 8.925 1.04 ;
      RECT 6.705 1.26 7.935 1.43 ;
      RECT 6.705 0.84 7.035 1.26 ;
      RECT 7.685 0.425 7.935 1.26 ;
      RECT 2.235 2.43 7.15 2.53 ;
      RECT 6.87 2.53 7.15 2.735 ;
      RECT 0.89 2.36 7.15 2.43 ;
      RECT 6.82 2.11 7.15 2.36 ;
      RECT 6.82 1.94 8.38 2.11 ;
      RECT 8.01 2.11 8.38 2.735 ;
      RECT 2.235 2.53 2.565 2.9 ;
      RECT 0.89 2.43 1.22 2.9 ;
      RECT 0.89 2.26 2.565 2.36 ;
      RECT 5.47 2.905 8.83 3.075 ;
      RECT 5.47 2.7 6.7 2.905 ;
      RECT 7.425 2.28 7.755 2.905 ;
      RECT 8.58 1.94 8.83 2.905 ;
      RECT 2.85 2.09 4.525 2.19 ;
      RECT 0.125 1.92 4.525 2.09 ;
      RECT 0.125 1.18 0.355 1.92 ;
      RECT 5.92 1.6 8.445 1.77 ;
      RECT 8.115 0.595 8.445 1.6 ;
      RECT 5.92 1.77 6.25 2.19 ;
      RECT 5.92 1.3 6.09 1.6 ;
      RECT 4.71 1.13 6.09 1.3 ;
      RECT 5.61 0.58 5.94 1.13 ;
      RECT 4.71 1.3 4.88 1.35 ;
      RECT 3.595 1.35 4.88 1.58 ;
      RECT 0.745 1.58 4.88 1.75 ;
      RECT 0.745 1.075 1.075 1.58 ;
      RECT 3.005 1.18 3.235 1.41 ;
      RECT 3.005 1.01 4.54 1.18 ;
      RECT 4.29 0.48 4.54 1.01 ;
      RECT 3.43 0.44 3.76 1.01 ;
      RECT 0 -0.085 9.6 0.085 ;
      RECT 7.215 0.085 7.465 1.09 ;
      RECT 6.13 0.085 6.3 0.675 ;
      RECT 3 0.085 3.25 0.84 ;
      RECT 3.94 0.085 4.11 0.84 ;
      RECT 4.72 0.085 5.44 0.96 ;
      RECT 6.275 0.96 6.525 1.28 ;
      RECT 6.13 0.675 6.525 0.96 ;
      RECT 1.935 0.085 2.105 0.675 ;
      RECT 1.935 0.675 2.33 1.07 ;
      RECT 0 3.245 9.6 3.415 ;
      RECT 2.845 2.7 3.175 3.245 ;
      RECT 3.745 2.7 4.075 3.245 ;
      RECT 4.645 2.7 4.975 3.245 ;
      RECT 1.395 2.6 2.065 3.245 ;
      RECT 0.32 2.26 0.65 3.245 ;
    LAYER mcon ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 1.21 0.325 1.38 ;
      RECT 3.035 1.21 3.205 1.38 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
  END
END scs8ls_a221o_4

MACRO scs8ls_a221oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.18 3.715 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505 1.35 2.835 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965 1.35 2.295 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.35 1.795 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.35 1.09 1.01 ;
        RECT 0.125 1.01 2.575 1.18 ;
        RECT 0.125 1.18 0.375 2.98 ;
        RECT 2.16 0.35 2.575 1.01 ;
    END
    ANTENNADIFFAREA 1.1775 ;
  END Y

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.35 0.875 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END C1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.275 2.12 1.545 2.735 ;
      RECT 1.275 1.95 3.525 2.12 ;
      RECT 2.255 2.12 2.505 2.98 ;
      RECT 3.195 2.12 3.525 2.98 ;
      RECT 3.195 1.82 3.525 1.95 ;
      RECT 0.575 2.905 2.055 3.075 ;
      RECT 1.725 2.29 2.055 2.905 ;
      RECT 0.575 1.95 0.905 2.905 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 3.17 0.085 3.5 1.01 ;
      RECT 1.26 0.085 1.63 0.825 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 2.675 2.29 3.025 3.245 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a221oi_1

MACRO scs8ls_a221oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585 1.35 0.915 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END C1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.895 1.43 5.635 1.78 ;
        RECT 4.895 1.78 5.065 1.95 ;
        RECT 3.405 1.95 5.065 2.12 ;
        RECT 3.405 1.43 3.735 1.95 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.43 4.675 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.55 3.235 1.95 ;
        RECT 1.425 1.95 3.235 2.12 ;
        RECT 2.685 1.43 3.015 1.55 ;
        RECT 1.425 1.68 1.595 1.95 ;
        RECT 1.245 1.43 1.595 1.68 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945 1.43 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.38 1.95 ;
        RECT 0.125 1.95 0.885 2.12 ;
        RECT 0.125 1.09 5.43 1.18 ;
        RECT 0.555 2.12 0.885 2.735 ;
        RECT 1.09 1.18 5.43 1.26 ;
        RECT 0.125 1.01 1.26 1.09 ;
        RECT 2.95 0.35 3.18 1.09 ;
        RECT 5.18 0.35 5.43 1.09 ;
        RECT 0.125 0.35 0.38 1.01 ;
        RECT 1.09 0.35 1.26 1.01 ;
    END
    ANTENNADIFFAREA 1.1722 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 0.56 0.085 0.91 0.84 ;
      RECT 1.94 0.085 2.28 0.58 ;
      RECT 4.2 0.085 4.53 0.58 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 3.355 2.63 3.605 3.245 ;
      RECT 4.335 2.63 4.505 3.245 ;
      RECT 5.235 1.95 5.485 3.245 ;
      RECT 3.35 0.75 5 0.92 ;
      RECT 3.35 0.33 4.03 0.75 ;
      RECT 4.7 0.33 5 0.75 ;
      RECT 1.44 0.75 2.78 0.92 ;
      RECT 1.44 0.35 1.77 0.75 ;
      RECT 2.45 0.33 2.78 0.75 ;
      RECT 1.455 2.46 1.815 2.735 ;
      RECT 1.455 2.29 5.035 2.46 ;
      RECT 3.805 2.46 4.135 2.98 ;
      RECT 4.705 2.46 5.035 2.98 ;
      RECT 0.105 2.905 3.165 2.98 ;
      RECT 2.015 2.63 3.165 2.905 ;
      RECT 1.085 1.85 1.255 2.905 ;
      RECT 0.105 2.98 2.265 3.075 ;
      RECT 0.105 2.29 0.355 2.905 ;
    LAYER mcon ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a221oi_2

MACRO scs8ls_a221oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.43 6.115 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.43 4.265 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.43 8.095 1.78 ;
        RECT 6.73 1.35 8.095 1.43 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285 1.35 9.955 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.35 1.875 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END C1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.35 0.495 1.01 ;
        RECT 0.105 1.01 2.295 1.09 ;
        RECT 0.105 1.09 8.21 1.18 ;
        RECT 1.185 0.35 1.355 1.01 ;
        RECT 2.045 0.35 2.295 1.01 ;
        RECT 0.105 1.18 0.355 2.905 ;
        RECT 2.045 1.18 6.53 1.26 ;
        RECT 6.36 0.85 8.21 1.09 ;
        RECT 4.85 0.64 5.04 1.09 ;
        RECT 5.71 0.64 5.9 1.09 ;
        RECT 0.105 2.905 2.235 3.075 ;
        RECT 7.915 0.77 8.21 0.85 ;
        RECT 1.005 2.29 1.335 2.905 ;
        RECT 1.905 2.29 2.235 2.905 ;
    END
    ANTENNADIFFAREA 2.3802 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 4.43 0.3 6.4 0.47 ;
      RECT 6.07 0.47 6.4 0.68 ;
      RECT 2.63 0.75 4.68 0.92 ;
      RECT 4.43 0.47 4.68 0.75 ;
      RECT 2.63 0.35 2.88 0.75 ;
      RECT 3.57 0.35 3.74 0.75 ;
      RECT 5.21 0.47 5.54 0.92 ;
      RECT 8.39 1.01 10.36 1.18 ;
      RECT 8.39 0.6 8.56 1.01 ;
      RECT 9.25 0.35 9.42 1.01 ;
      RECT 10.11 0.35 10.36 1.01 ;
      RECT 6.59 0.35 8.56 0.6 ;
      RECT 6.59 0.6 6.92 0.68 ;
      RECT 7.45 0.6 7.745 0.68 ;
      RECT 2.615 2.46 2.945 2.98 ;
      RECT 2.615 2.29 6.725 2.46 ;
      RECT 3.515 2.46 3.845 2.98 ;
      RECT 4.415 2.46 4.745 2.98 ;
      RECT 5.315 2.46 5.645 2.98 ;
      RECT 6.445 2.46 6.725 2.905 ;
      RECT 6.445 2.905 10.375 3.075 ;
      RECT 7.395 2.29 7.625 2.905 ;
      RECT 8.295 2.29 8.525 2.905 ;
      RECT 9.195 2.29 9.425 2.905 ;
      RECT 10.125 1.82 10.375 2.905 ;
      RECT 0.555 1.95 9.925 2.12 ;
      RECT 6.895 2.12 7.225 2.735 ;
      RECT 7.795 2.12 8.125 2.735 ;
      RECT 8.695 2.12 9.025 2.735 ;
      RECT 9.595 2.12 9.925 2.735 ;
      RECT 0.555 2.12 0.835 2.735 ;
      RECT 1.505 2.12 1.735 2.735 ;
      RECT 0 -0.085 10.56 0.085 ;
      RECT 8.74 0.085 9.07 0.84 ;
      RECT 9.6 0.085 9.93 0.84 ;
      RECT 0.675 0.085 1.005 0.84 ;
      RECT 1.535 0.085 1.865 0.84 ;
      RECT 3.06 0.085 3.39 0.58 ;
      RECT 3.92 0.085 4.25 0.58 ;
      RECT 0 3.245 10.56 3.415 ;
      RECT 3.145 2.63 3.315 3.245 ;
      RECT 4.045 2.63 4.215 3.245 ;
      RECT 4.945 2.63 5.115 3.245 ;
      RECT 5.815 2.63 6.275 3.245 ;
    LAYER mcon ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
  END
END scs8ls_a221oi_4

MACRO scs8ls_a222o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.22 1.12 2.755 1.79 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.12 3.255 1.52 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.12 3.825 1.545 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.18 1.93 1.76 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.12 0.55 1.79 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END C1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.355 1.82 4.71 2.98 ;
        RECT 4.54 1.13 4.71 1.82 ;
        RECT 4.355 0.35 4.71 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
  END X

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.06 1.12 1.39 1.76 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END C2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 0.96 0.085 1.805 0.6 ;
      RECT 3.62 0.085 4.185 0.61 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 2.82 2.3 3.15 3.245 ;
      RECT 3.855 1.895 4.185 3.245 ;
      RECT 1.72 2.13 2.05 2.735 ;
      RECT 1.72 1.96 3.65 2.13 ;
      RECT 3.32 2.13 3.65 2.935 ;
      RECT 1.72 1.93 2.05 1.96 ;
      RECT 3.32 1.895 3.65 1.96 ;
      RECT 0.115 2.905 2.59 3.075 ;
      RECT 2.26 2.3 2.59 2.905 ;
      RECT 0.115 1.96 0.445 2.905 ;
      RECT 1.22 1.93 1.55 2.905 ;
      RECT 4.015 1.3 4.37 1.63 ;
      RECT 0.14 0.78 4.185 0.95 ;
      RECT 4.015 0.95 4.185 1.3 ;
      RECT 2.295 0.33 3.13 0.78 ;
      RECT 0.72 1.93 1.05 2.735 ;
      RECT 0.72 0.95 0.89 1.93 ;
      RECT 0.14 0.35 0.47 0.78 ;
    LAYER mcon ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a222o_1

MACRO scs8ls_a222o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.35 3.255 2.15 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.26 1.14 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END C2

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.685 1.35 5.155 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.465 1.35 3.795 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.35 4.445 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.3 0.435 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END C1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 1.82 2.44 2.2 ;
        RECT 1.695 0.92 2.025 1.82 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.935 0.085 1.185 0.75 ;
      RECT 0 -0.085 5.28 0.085 ;
      RECT 2.205 0.085 2.535 0.41 ;
      RECT 4.26 0.085 4.59 0.84 ;
      RECT 0 3.245 5.28 3.415 ;
      RECT 2.645 2.71 2.975 3.245 ;
      RECT 4.835 1.95 5.165 3.245 ;
      RECT 1.575 2.71 1.905 3.245 ;
      RECT 3.265 2.905 4.665 3.075 ;
      RECT 3.265 2.71 3.63 2.905 ;
      RECT 4.335 1.95 4.665 2.905 ;
      RECT 0.565 2.37 4.165 2.54 ;
      RECT 3.835 2.54 4.165 2.735 ;
      RECT 3.835 1.95 4.165 2.37 ;
      RECT 0.565 2.54 0.895 2.98 ;
      RECT 2.23 1.01 3.75 1.18 ;
      RECT 3.265 0.7 3.75 1.01 ;
      RECT 1.355 0.58 2.4 0.75 ;
      RECT 2.23 0.75 2.4 1.01 ;
      RECT 2.23 1.18 2.56 1.59 ;
      RECT 0.115 1.95 1.525 2.2 ;
      RECT 1.355 1.09 1.525 1.95 ;
      RECT 0.115 0.92 1.525 1.09 ;
      RECT 1.355 0.75 1.525 0.92 ;
      RECT 0.115 2.2 0.365 2.98 ;
      RECT 0.115 0.39 0.365 0.92 ;
      RECT 3.92 1.01 5.14 1.18 ;
      RECT 3.92 0.52 4.09 1.01 ;
      RECT 4.81 0.35 5.14 1.01 ;
      RECT 2.765 0.35 4.09 0.52 ;
      RECT 2.765 0.52 3.095 0.84 ;
    LAYER mcon ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a222o_2

MACRO scs8ls_a222oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975 1.12 2.305 1.79 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.14 0.78 3.36 0.95 ;
        RECT 1.485 0.95 1.795 1.78 ;
        RECT 0.14 0.35 0.47 0.78 ;
        RECT 2.525 0.33 3.36 0.78 ;
        RECT 1.485 1.78 1.655 1.96 ;
        RECT 0.115 1.96 1.655 2.13 ;
        RECT 0.115 2.13 0.445 2.98 ;
        RECT 1.115 2.13 1.655 2.735 ;
    END
    ANTENNADIFFAREA 1.232 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.155 1.12 3.715 1.79 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885 1.18 4.215 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.12 2.875 1.79 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.12 0.595 1.79 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985 1.12 1.315 1.79 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END C2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.615 2.905 2.655 3.075 ;
      RECT 2.325 2.3 2.655 2.905 ;
      RECT 0.615 2.3 0.945 2.905 ;
      RECT 1.825 2.13 2.155 2.735 ;
      RECT 1.825 1.96 4.205 2.13 ;
      RECT 2.825 2.13 3.155 2.98 ;
      RECT 3.875 2.13 4.205 2.98 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 3.85 0.085 4.18 0.95 ;
      RECT 0.96 0.085 2.18 0.6 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 3.325 2.3 3.655 3.245 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a222oi_1

MACRO scs8ls_a222oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.675 1.47 3.235 1.8 ;
        RECT 3.065 1.8 3.235 1.95 ;
        RECT 3.065 1.95 4.275 2.12 ;
        RECT 4.105 1.78 4.275 1.95 ;
        RECT 4.105 1.45 4.475 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.165 0.835 1.495 ;
        RECT 0.605 1.495 0.835 1.665 ;
        RECT 0.605 1.665 2.125 1.835 ;
        RECT 1.795 1.13 2.125 1.665 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END C2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 2.005 2.465 2.175 ;
        RECT 0.085 2.175 0.365 2.98 ;
        RECT 1.065 2.175 1.325 2.735 ;
        RECT 1.995 2.175 2.465 2.735 ;
        RECT 0.085 1.92 0.365 2.005 ;
        RECT 2.295 1.3 2.465 2.005 ;
        RECT 0.085 0.995 0.255 1.92 ;
        RECT 2.295 1.13 2.84 1.3 ;
        RECT 0.085 0.825 1.42 0.995 ;
        RECT 2.51 1.09 2.84 1.13 ;
        RECT 1.09 0.78 1.42 0.825 ;
        RECT 2.51 0.92 4.715 1.09 ;
        RECT 4.45 1.09 4.715 1.11 ;
        RECT 2.51 0.35 2.84 0.92 ;
        RECT 4.45 0.35 4.715 0.92 ;
        RECT 4.45 1.11 6.58 1.28 ;
        RECT 6.32 0.35 6.58 1.11 ;
    END
    ANTENNADIFFAREA 1.6932 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.45 6.455 1.78 ;
        RECT 5.885 1.78 6.055 1.95 ;
        RECT 4.945 1.95 6.055 2.12 ;
        RECT 4.945 1.78 5.115 1.95 ;
        RECT 4.685 1.45 5.115 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.305 1.45 5.635 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.26 3.735 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.165 1.335 1.495 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END C1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.72 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.72 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.02 0.58 4.27 0.75 ;
      RECT 3.02 0.35 3.27 0.58 ;
      RECT 4.02 0.35 4.27 0.58 ;
      RECT 4.885 0.77 6.15 0.94 ;
      RECT 4.885 0.35 5.215 0.77 ;
      RECT 5.9 0.33 6.15 0.77 ;
      RECT 1.59 0.61 1.78 0.885 ;
      RECT 0.66 0.35 1.78 0.61 ;
      RECT 0.565 2.98 3.335 3.075 ;
      RECT 0.565 2.905 4.325 2.98 ;
      RECT 3.005 2.65 4.325 2.905 ;
      RECT 3.005 2.63 3.335 2.65 ;
      RECT 0.565 2.345 0.895 2.905 ;
      RECT 1.495 2.345 1.825 2.905 ;
      RECT 4.5 2.46 6.605 2.48 ;
      RECT 5.425 2.48 5.655 2.98 ;
      RECT 6.335 2.48 6.605 3 ;
      RECT 2.635 2.29 6.605 2.46 ;
      RECT 6.275 1.95 6.605 2.29 ;
      RECT 4.5 2.48 4.715 2.98 ;
      RECT 4.445 1.95 4.775 2.29 ;
      RECT 2.635 2.46 2.805 2.735 ;
      RECT 2.635 1.97 2.805 2.29 ;
      RECT 0 -0.085 6.72 0.085 ;
      RECT 0.115 0.085 0.48 0.655 ;
      RECT 1.95 0.085 2.28 0.94 ;
      RECT 3.45 0.085 3.84 0.41 ;
      RECT 5.385 0.085 5.715 0.6 ;
      RECT 0 3.245 6.72 3.415 ;
      RECT 4.895 2.65 5.255 3.245 ;
      RECT 5.825 2.65 6.155 3.245 ;
    LAYER mcon ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a222oi_2

MACRO scs8ls_a22o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965 1.35 2.295 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.505 0.355 0.67 ;
        RECT 0.125 0.255 0.56 0.505 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.425 1.47 1.795 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.47 1.215 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B2

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 0.35 3.255 2.98 ;
    END
    ANTENNADIFFAREA 0.5041 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.645 2.905 1.995 3.075 ;
      RECT 1.595 2.31 1.995 2.905 ;
      RECT 0.645 1.97 0.895 2.905 ;
      RECT 0.22 1.13 1.285 1.3 ;
      RECT 0.22 0.84 0.55 1.13 ;
      RECT 1.115 0.625 1.285 1.13 ;
      RECT 1.115 0.375 2.245 0.625 ;
      RECT 1.095 1.97 2.755 2.14 ;
      RECT 2.505 1.18 2.755 1.97 ;
      RECT 1.485 1.01 2.755 1.18 ;
      RECT 1.095 2.14 1.425 2.735 ;
      RECT 1.485 0.795 1.815 1.01 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 0.73 0.085 0.945 0.96 ;
      RECT 2.495 0.085 2.745 0.84 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.165 2.31 2.725 3.245 ;
      RECT 0.195 1.97 0.445 3.245 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a22o_1

MACRO scs8ls_a22o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585 1.35 1.905 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.35 3.735 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075 1.35 2.495 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.705 1.35 3.235 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B2

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.53 0.35 0.86 1.72 ;
        RECT 0.53 1.72 1.075 1.89 ;
        RECT 0.905 1.89 1.075 2.29 ;
        RECT 0.905 2.29 1.185 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.925 2.905 3.225 3.075 ;
      RECT 1.925 2.29 2.255 2.905 ;
      RECT 2.875 1.95 3.225 2.905 ;
      RECT 2.5 1.01 3.7 1.18 ;
      RECT 2.5 0.425 2.67 1.01 ;
      RECT 3.37 0.35 3.7 1.01 ;
      RECT 1.5 0.255 2.67 0.425 ;
      RECT 1.5 0.425 1.83 0.84 ;
      RECT 2.455 2.12 2.705 2.735 ;
      RECT 1.245 1.95 2.705 2.12 ;
      RECT 1.085 1.01 2.33 1.18 ;
      RECT 2 0.595 2.33 1.01 ;
      RECT 1.245 1.55 1.415 1.95 ;
      RECT 1.085 1.18 1.415 1.55 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 1.04 0.085 1.29 0.84 ;
      RECT 2.87 0.085 3.2 0.84 ;
      RECT 0.1 0.085 0.35 1.13 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 1.385 2.29 1.715 3.245 ;
      RECT 3.395 1.95 3.725 3.245 ;
      RECT 0.485 2.06 0.735 3.245 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a22o_2

MACRO scs8ls_a22o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405 1.45 6.115 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.955 0.255 5.32 0.505 ;
        RECT 4.955 0.505 5.125 0.67 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.495 1.435 3.825 1.765 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.155 1.935 4.195 2.15 ;
        RECT 4.025 1.77 4.195 1.935 ;
        RECT 3.155 1.765 3.325 1.935 ;
        RECT 4.025 1.44 4.655 1.77 ;
        RECT 3.025 1.435 3.325 1.765 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B2

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 1.855 1.41 ;
        RECT 0.705 1.41 1.855 1.65 ;
        RECT 0.125 1.14 2.515 1.18 ;
        RECT 0.705 1.65 0.875 2.98 ;
        RECT 1.525 1.65 1.855 2.98 ;
        RECT 1.405 1.01 2.515 1.14 ;
        RECT 1.405 0.48 1.655 1.01 ;
        RECT 2.265 0.48 2.515 1.01 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 4.14 0.83 4.355 0.925 ;
      RECT 3.2 0.58 4.355 0.83 ;
      RECT 2.815 2.32 4.865 2.49 ;
      RECT 4.615 2.49 4.865 2.98 ;
      RECT 4.615 2.12 4.865 2.32 ;
      RECT 4.615 1.95 6.91 2.12 ;
      RECT 5.68 2.12 5.93 2.98 ;
      RECT 6.66 2.12 6.91 2.98 ;
      RECT 4.615 1.94 4.865 1.95 ;
      RECT 6.66 1.94 6.91 1.95 ;
      RECT 2.815 2.49 2.985 2.735 ;
      RECT 2.815 1.94 2.985 2.32 ;
      RECT 2.685 1.095 6.055 1.265 ;
      RECT 5.725 1.265 6.055 1.275 ;
      RECT 5.725 1.015 6.055 1.095 ;
      RECT 2.475 2.905 4.415 2.98 ;
      RECT 3.185 2.66 4.415 2.905 ;
      RECT 2.475 1.68 2.645 2.905 ;
      RECT 2.025 1.35 2.855 1.68 ;
      RECT 2.685 1.265 2.855 1.35 ;
      RECT 2.475 2.98 3.515 3.075 ;
      RECT 3.63 1 3.96 1.095 ;
      RECT 0 -0.085 7.2 0.085 ;
      RECT 6.585 0.085 6.915 1.275 ;
      RECT 2.695 0.085 3.025 0.925 ;
      RECT 4.535 0.085 4.785 0.925 ;
      RECT 0.975 0.085 1.225 0.97 ;
      RECT 1.835 0.085 2.085 0.84 ;
      RECT 0 3.245 7.2 3.415 ;
      RECT 5.035 2.29 5.51 3.245 ;
      RECT 6.13 2.29 6.46 3.245 ;
      RECT 2.055 1.85 2.305 3.245 ;
      RECT 0.175 1.9 0.505 3.245 ;
      RECT 1.075 1.82 1.325 3.245 ;
      RECT 6.235 0.845 6.405 1.275 ;
      RECT 5.295 0.675 6.405 0.845 ;
      RECT 6.235 0.595 6.405 0.675 ;
    LAYER mcon ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a22o_4

MACRO scs8ls_a22oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.35 1.875 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.35 1.335 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.18 0.835 1.95 ;
        RECT 0.605 1.95 1.015 2.12 ;
        RECT 0.605 1.01 1.57 1.18 ;
        RECT 0.845 2.12 1.015 2.735 ;
        RECT 1.13 0.35 1.57 1.01 ;
    END
    ANTENNADIFFAREA 0.6246 ;
  END Y

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.435 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.315 2.905 1.545 3.075 ;
      RECT 1.215 2.12 1.545 2.905 ;
      RECT 1.215 1.95 2.565 2.12 ;
      RECT 2.235 2.12 2.565 2.98 ;
      RECT 0.315 2.29 0.645 2.905 ;
      RECT 0 -0.085 2.88 0.085 ;
      RECT 2.21 0.085 2.54 1.13 ;
      RECT 0.34 0.085 0.67 0.84 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 1.715 2.29 2.065 3.245 ;
    LAYER mcon ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a22oi_1

MACRO scs8ls_a22oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.72 1.26 3.235 1.55 ;
        RECT 2.72 1.09 4.075 1.26 ;
        RECT 3.905 1.26 4.075 1.3 ;
        RECT 3.905 1.3 4.37 1.63 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.04 0.81 2.55 1.09 ;
        RECT 0.285 1.09 2.55 1.26 ;
        RECT 2.145 0.35 2.55 0.81 ;
        RECT 2.38 1.26 2.55 1.72 ;
        RECT 0.285 0.35 0.535 1.09 ;
        RECT 2.38 1.72 3.13 1.89 ;
        RECT 2.93 1.89 3.13 1.95 ;
        RECT 2.93 1.95 4.71 2.12 ;
        RECT 2.93 2.12 3.13 2.735 ;
        RECT 3.86 2.12 4.03 2.735 ;
        RECT 4.54 1.13 4.71 1.95 ;
        RECT 4.245 0.35 4.71 1.13 ;
    END
    ANTENNADIFFAREA 1.4974 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.43 0.88 1.78 ;
        RECT 0.71 1.78 0.88 1.95 ;
        RECT 0.71 1.95 2.21 2.12 ;
        RECT 1.88 1.43 2.21 1.95 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.05 1.43 1.42 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.43 3.735 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.835 0.75 4.065 0.92 ;
      RECT 2.835 0.33 3.135 0.75 ;
      RECT 3.815 0.33 4.065 0.75 ;
      RECT 2.4 2.905 4.56 3.075 ;
      RECT 4.23 2.29 4.56 2.905 ;
      RECT 0.29 2.29 2.73 2.46 ;
      RECT 1.19 2.46 1.52 2.98 ;
      RECT 2.4 2.46 2.73 2.905 ;
      RECT 2.4 2.06 2.73 2.29 ;
      RECT 3.33 2.29 3.66 2.905 ;
      RECT 0.29 2.46 0.54 2.98 ;
      RECT 0.29 1.95 0.54 2.29 ;
      RECT 0.715 0.75 1.815 0.92 ;
      RECT 1.645 0.64 1.815 0.75 ;
      RECT 0.715 0.33 0.965 0.75 ;
      RECT 1.645 0.35 1.975 0.64 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 1.145 0.085 1.475 0.58 ;
      RECT 3.305 0.085 3.635 0.58 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 0.74 2.63 0.99 3.245 ;
      RECT 1.69 2.63 2.23 3.245 ;
    LAYER mcon ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a22oi_2

MACRO scs8ls_a22oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.35 5.635 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.35 7.465 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.265 1.35 3.275 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.35 1.955 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.445 1.18 4.195 1.52 ;
        RECT 3.445 1.52 3.615 1.95 ;
        RECT 2.35 1.13 4.195 1.18 ;
        RECT 0.635 1.95 3.615 2.12 ;
        RECT 2.35 1.01 5.78 1.13 ;
        RECT 0.635 2.12 0.885 2.735 ;
        RECT 1.615 2.12 1.785 2.735 ;
        RECT 2.515 2.12 2.685 2.735 ;
        RECT 3.415 2.12 3.615 2.735 ;
        RECT 3.21 0.85 5.78 1.01 ;
        RECT 2.35 0.595 2.68 1.01 ;
        RECT 3.21 0.77 3.99 0.85 ;
        RECT 5.45 0.77 5.78 0.85 ;
    END
    ANTENNADIFFAREA 2.1728 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 5.96 1.01 7.93 1.18 ;
      RECT 5.96 0.6 6.13 1.01 ;
      RECT 6.74 0.35 6.99 1.01 ;
      RECT 7.6 0.35 7.93 1.01 ;
      RECT 4.16 0.35 6.13 0.6 ;
      RECT 4.16 0.6 4.49 0.68 ;
      RECT 2 0.255 3.97 0.425 ;
      RECT 2.86 0.425 3.97 0.6 ;
      RECT 0.2 1.01 2.17 1.18 ;
      RECT 2 0.425 2.17 1.01 ;
      RECT 0.2 0.35 0.45 1.01 ;
      RECT 1.06 0.35 1.31 1.01 ;
      RECT 2.86 0.6 3.03 0.84 ;
      RECT 0.185 2.905 4.035 3.075 ;
      RECT 3.785 2.12 4.035 2.905 ;
      RECT 3.785 1.95 7.945 2.12 ;
      RECT 4.765 2.12 5.015 2.98 ;
      RECT 5.815 2.12 6.065 2.98 ;
      RECT 6.795 2.12 6.965 2.98 ;
      RECT 7.695 2.12 7.945 2.98 ;
      RECT 3.785 1.82 4.035 1.95 ;
      RECT 7.695 1.82 7.945 1.95 ;
      RECT 0.185 1.82 0.435 2.905 ;
      RECT 1.085 2.29 1.415 2.905 ;
      RECT 1.985 2.29 2.315 2.905 ;
      RECT 2.885 2.29 3.215 2.905 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 6.31 0.085 6.56 0.84 ;
      RECT 7.17 0.085 7.42 0.84 ;
      RECT 0.63 0.085 0.88 0.84 ;
      RECT 1.49 0.085 1.82 0.84 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 4.235 2.29 4.565 3.245 ;
      RECT 5.185 2.29 5.645 3.245 ;
      RECT 6.265 2.29 6.595 3.245 ;
      RECT 7.165 2.29 7.495 3.245 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
  END
END scs8ls_a22oi_4

MACRO scs8ls_a2bb2o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.18 1.85 1.62 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END A2N

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 0.255 4.195 0.67 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.82 0.56 2.98 ;
        RECT 0.125 1.15 0.295 1.82 ;
        RECT 0.125 0.42 0.59 1.15 ;
    END
    ANTENNADIFFAREA 0.5041 ;
  END X

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 1.18 1.335 1.62 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END A1N

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.875 1.45 3.235 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.715 2.12 2.885 2.98 ;
      RECT 2.715 1.95 3.895 2.12 ;
      RECT 3.645 2.12 3.895 2.98 ;
      RECT 3.645 1.94 3.895 1.95 ;
      RECT 1.285 0.52 1.59 1.01 ;
      RECT 1.285 0.255 2.595 0.52 ;
      RECT 2.02 1.03 2.9 1.21 ;
      RECT 1.325 2.905 2.515 3.075 ;
      RECT 2.185 2.47 2.515 2.905 ;
      RECT 0.73 1.79 2.19 1.96 ;
      RECT 2.02 1.21 2.19 1.79 ;
      RECT 1.325 1.96 1.495 2.905 ;
      RECT 0.73 1.65 0.9 1.79 ;
      RECT 0.465 1.32 0.9 1.65 ;
      RECT 1.665 2.3 1.995 2.735 ;
      RECT 1.665 2.13 2.53 2.3 ;
      RECT 2.36 1.78 2.53 2.13 ;
      RECT 2.36 1.45 2.665 1.78 ;
      RECT 3.54 1.01 3.87 1.29 ;
      RECT 3.145 0.84 3.87 1.01 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 3.145 0.085 3.315 0.84 ;
      RECT 2.765 0.085 2.935 0.69 ;
      RECT 1.76 0.69 2.935 0.86 ;
      RECT 0.77 0.085 1.1 1.01 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 3.085 2.29 3.445 3.245 ;
      RECT 0.76 2.13 1.09 3.245 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a2bb2o_1

MACRO scs8ls_a2bb2o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.18 3.255 2.15 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END A1N

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 0.35 3.92 2.15 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.385 1.18 2.755 1.51 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END A2N

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.435 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.18 1.315 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 3.105 2.66 3.495 3.245 ;
      RECT 4.065 2.66 4.395 3.245 ;
      RECT 0.715 2.06 1.045 3.245 ;
      RECT 0.265 1.89 0.515 2.98 ;
      RECT 0.265 1.72 1.415 1.89 ;
      RECT 1.245 1.89 1.415 2.98 ;
      RECT 2.265 1.85 2.58 2.64 ;
      RECT 1.925 1.68 2.58 1.85 ;
      RECT 1.925 0.84 2.87 1.01 ;
      RECT 2.69 0.35 2.87 0.84 ;
      RECT 1.925 1.01 2.175 1.68 ;
      RECT 2.75 2.32 4.47 2.49 ;
      RECT 4.09 1.35 4.47 2.32 ;
      RECT 1.585 2.81 2.92 2.98 ;
      RECT 2.75 2.49 2.92 2.81 ;
      RECT 1.585 2.02 1.945 2.81 ;
      RECT 1.585 1.55 1.755 2.02 ;
      RECT 1.485 1.38 1.755 1.55 ;
      RECT 1.485 1.01 1.655 1.38 ;
      RECT 1.08 0.84 1.655 1.01 ;
      RECT 1.08 0.35 1.48 0.84 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 4.1 0.085 4.35 1.13 ;
      RECT 0.29 0.085 0.62 1.01 ;
      RECT 1.65 0.085 2.52 0.67 ;
      RECT 3.05 0.085 3.315 0.94 ;
    LAYER mcon ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a2bb2o_2

MACRO scs8ls_a2bb2o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555 1.35 2.85 1.78 ;
    END
    ANTENNAGATEAREA 0.264 ;
  END A1N

  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.36 1.35 3.685 1.78 ;
    END
    ANTENNAGATEAREA 0.264 ;
  END A2N

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.26 7.075 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405 1.26 6.115 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B2

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.13 0.835 1.78 ;
        RECT 0.665 1.78 0.835 1.8 ;
        RECT 0.125 0.96 2.045 1.13 ;
        RECT 0.665 1.8 2.24 1.97 ;
        RECT 0.935 0.35 1.185 0.96 ;
        RECT 1.795 0.35 2.045 0.96 ;
        RECT 1.01 1.97 1.34 2.98 ;
        RECT 1.91 1.97 2.24 2.98 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 4.06 2.905 5.21 3.075 ;
      RECT 4.06 2.29 4.39 2.905 ;
      RECT 4.96 2.12 5.21 2.905 ;
      RECT 4.96 1.95 7.09 2.12 ;
      RECT 5.86 2.12 6.19 2.98 ;
      RECT 6.76 2.12 7.09 2.98 ;
      RECT 3.29 2.12 3.62 2.98 ;
      RECT 3.02 1.95 4.15 2.12 ;
      RECT 3.855 1.47 4.15 1.95 ;
      RECT 3.02 1.13 3.19 1.95 ;
      RECT 2.985 0.595 3.19 1.13 ;
      RECT 4.565 0.35 5.765 0.6 ;
      RECT 2.645 0.255 3.53 0.425 ;
      RECT 3.36 0.425 3.53 1.01 ;
      RECT 3.36 1.01 4.815 1.18 ;
      RECT 4.565 1.18 4.76 2.735 ;
      RECT 4.565 0.6 4.815 1.01 ;
      RECT 2.215 1.01 2.815 1.18 ;
      RECT 2.645 0.425 2.815 1.01 ;
      RECT 1.035 1.3 2.385 1.63 ;
      RECT 2.215 1.18 2.385 1.3 ;
      RECT 6.295 0.35 6.665 0.75 ;
      RECT 6.495 0.085 6.665 0.35 ;
      RECT 0 -0.085 7.2 0.085 ;
      RECT 2.225 0.085 2.475 0.84 ;
      RECT 3.7 0.085 4.385 0.84 ;
      RECT 0.505 0.085 0.755 0.79 ;
      RECT 1.365 0.085 1.615 0.79 ;
      RECT 0 3.245 7.2 3.415 ;
      RECT 5.41 2.29 5.66 3.245 ;
      RECT 6.39 2.29 6.56 3.245 ;
      RECT 2.41 1.95 2.78 3.245 ;
      RECT 0.56 2.14 0.81 3.245 ;
      RECT 1.54 2.14 1.71 3.245 ;
      RECT 5.005 0.92 7.095 1.09 ;
      RECT 5.005 0.77 6.115 0.92 ;
      RECT 6.845 0.35 7.095 0.92 ;
      RECT 5.945 0.35 6.115 0.77 ;
    LAYER mcon ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a2bb2o_4

MACRO scs8ls_a2bb2oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.18 3.255 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.54 2.755 2.15 ;
        RECT 2.22 1.22 2.755 1.54 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B2

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.26 0.435 1.78 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END A1N

  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.45 1.1 1.78 ;
    END
    ANTENNAGATEAREA 0.233 ;
  END A2N

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.61 1.92 2.275 2.22 ;
        RECT 1.61 2.22 1.78 2.29 ;
        RECT 1.61 1.75 2.05 1.92 ;
        RECT 1.53 2.29 1.78 2.98 ;
        RECT 1.88 1.05 2.05 1.75 ;
        RECT 1.88 0.88 2.315 1.05 ;
        RECT 2.055 0.35 2.315 0.88 ;
    END
    ANTENNADIFFAREA 0.5152 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.885 0.085 3.215 1.01 ;
      RECT 1.105 0.71 1.71 0.79 ;
      RECT 0.175 0.085 0.425 1.09 ;
      RECT 1.105 0.085 1.885 0.71 ;
      RECT 1.98 2.39 3.24 2.56 ;
      RECT 2.99 2.56 3.24 2.98 ;
      RECT 2.99 1.82 3.24 2.39 ;
      RECT 1.98 2.56 2.23 2.98 ;
      RECT 1.27 1.22 1.71 1.55 ;
      RECT 0.96 2.12 1.29 2.98 ;
      RECT 0.96 1.95 1.44 2.12 ;
      RECT 1.27 1.55 1.44 1.95 ;
      RECT 1.27 1.13 1.44 1.22 ;
      RECT 0.605 0.96 1.44 1.13 ;
      RECT 0.605 0.54 0.935 0.96 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.43 2.98 2.6 3.245 ;
      RECT 2.43 2.73 2.79 2.98 ;
      RECT 0.12 1.95 0.45 3.245 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a2bb2oi_1

MACRO scs8ls_a2bb2oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.285 0.435 0.67 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1N

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.35 4.675 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.32 3.735 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END B2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.15 3.235 1.41 ;
        RECT 2.525 1.41 2.78 2.735 ;
        RECT 2.08 0.98 3.795 1.15 ;
        RECT 3.465 0.77 3.795 0.98 ;
        RECT 2.08 0.39 2.25 0.98 ;
    END
    ANTENNADIFFAREA 0.7504 ;
  END Y

  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.45 1.57 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2N

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.08 2.905 3.23 3.075 ;
      RECT 2.98 2.12 3.23 2.905 ;
      RECT 2.98 1.95 5.11 2.12 ;
      RECT 3.96 2.12 4.13 2.98 ;
      RECT 4.86 2.12 5.11 2.98 ;
      RECT 2.98 1.82 3.23 1.95 ;
      RECT 4.86 1.82 5.11 1.95 ;
      RECT 2.08 1.82 2.33 2.905 ;
      RECT 3.975 1.01 5.085 1.18 ;
      RECT 3.975 0.6 4.145 1.01 ;
      RECT 4.755 0.35 5.085 1.01 ;
      RECT 3.035 0.35 4.145 0.6 ;
      RECT 1.74 1.32 2.205 1.65 ;
      RECT 1.42 1.95 1.91 2.98 ;
      RECT 1.74 1.65 1.91 1.95 ;
      RECT 1.74 1.28 1.91 1.32 ;
      RECT 1.035 1.11 1.91 1.28 ;
      RECT 1.035 0.49 1.33 1.11 ;
      RECT 0 -0.085 5.28 0.085 ;
      RECT 4.325 0.085 4.575 0.84 ;
      RECT 0.605 0.085 0.855 1.17 ;
      RECT 1.57 0.085 1.9 0.94 ;
      RECT 2.43 0.085 2.76 0.81 ;
      RECT 0 3.245 5.28 3.415 ;
      RECT 3.43 2.29 3.76 3.245 ;
      RECT 4.33 2.29 4.66 3.245 ;
      RECT 0.58 1.94 0.91 3.245 ;
    LAYER mcon ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a2bb2oi_2

MACRO scs8ls_a2bb2oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.47 2.275 1.8 ;
    END
    ANTENNAGATEAREA 0.411 ;
  END A1N

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.735 1.35 8.515 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.35 6.115 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END B2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.27 0.79 6.15 0.96 ;
        RECT 3.965 0.96 6.15 1.13 ;
        RECT 4.96 0.77 6.15 0.79 ;
        RECT 2.27 0.35 2.52 0.79 ;
        RECT 3.21 0.35 3.38 0.79 ;
        RECT 3.965 1.13 4.255 1.72 ;
        RECT 3.185 1.72 4.255 1.89 ;
        RECT 3.185 1.89 3.355 2.735 ;
        RECT 4.085 1.89 4.255 2.735 ;
    END
    ANTENNADIFFAREA 1.5008 ;
  END Y

  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.42 0.455 1.77 ;
    END
    ANTENNAGATEAREA 0.411 ;
  END A2N

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.105 2.905 1.255 3.075 ;
      RECT 1.085 2.14 1.255 2.905 ;
      RECT 0.105 1.94 0.435 2.905 ;
      RECT 1.085 1.97 2.235 2.14 ;
      RECT 1.905 2.14 2.235 2.98 ;
      RECT 1.085 1.94 1.255 1.97 ;
      RECT 2.655 2.905 4.785 3.075 ;
      RECT 4.455 2.12 4.785 2.905 ;
      RECT 4.455 1.95 8.385 2.12 ;
      RECT 5.355 2.12 5.685 2.98 ;
      RECT 6.335 2.12 6.505 2.98 ;
      RECT 7.155 2.12 7.485 2.98 ;
      RECT 8.055 2.12 8.385 2.98 ;
      RECT 6.335 1.82 6.505 1.95 ;
      RECT 2.655 1.82 2.985 2.905 ;
      RECT 3.555 2.06 3.885 2.905 ;
      RECT 0.635 1.13 3.585 1.3 ;
      RECT 2.575 1.3 3.585 1.55 ;
      RECT 1.45 0.35 1.62 1.13 ;
      RECT 0.635 1.3 0.885 2.735 ;
      RECT 6.33 1.01 8.3 1.18 ;
      RECT 6.33 0.6 6.5 1.01 ;
      RECT 7.11 0.35 7.36 1.01 ;
      RECT 7.97 0.35 8.3 1.01 ;
      RECT 4.53 0.35 6.5 0.6 ;
      RECT 0 -0.085 8.64 0.085 ;
      RECT 6.68 0.085 6.93 0.84 ;
      RECT 7.54 0.085 7.79 0.84 ;
      RECT 0.94 0.085 1.27 0.96 ;
      RECT 1.8 0.085 2.09 0.885 ;
      RECT 2.7 0.085 3.03 0.62 ;
      RECT 3.56 0.085 3.89 0.62 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 4.985 2.29 5.155 3.245 ;
      RECT 5.885 2.29 6.135 3.245 ;
      RECT 6.705 2.29 6.955 3.245 ;
      RECT 7.685 2.29 7.855 3.245 ;
      RECT 1.455 2.31 1.705 3.245 ;
    LAYER mcon ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
  END
END scs8ls_a2bb2oi_4

MACRO scs8ls_a311o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.44 2.335 0.67 ;
        RECT 2.005 0.255 2.335 0.44 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.45 1.905 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115 1.45 1.365 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 0.505 2.725 0.67 ;
        RECT 2.525 0.255 2.875 0.505 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385 0.255 3.715 0.67 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END C1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.85 0.475 2.98 ;
        RECT 0.125 1.18 0.295 1.85 ;
        RECT 0.125 1.01 0.605 1.18 ;
        RECT 0.355 0.48 0.605 1.01 ;
    END
    ANTENNADIFFAREA 0.5041 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.275 2.12 1.605 2.98 ;
      RECT 1.275 1.95 2.595 2.12 ;
      RECT 2.265 2.12 2.595 2.98 ;
      RECT 2.265 1.94 2.595 1.95 ;
      RECT 3.105 1.94 3.575 2.98 ;
      RECT 3.245 1.615 3.575 1.94 ;
      RECT 2.24 1.445 3.575 1.615 ;
      RECT 2.24 1.28 2.57 1.445 ;
      RECT 3.245 1.015 3.575 1.445 ;
      RECT 0.775 1.11 2.57 1.28 ;
      RECT 2.24 0.84 2.57 1.11 ;
      RECT 0.775 1.28 0.945 1.35 ;
      RECT 0.48 1.35 0.945 1.68 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 2.75 0.855 3.075 1.185 ;
      RECT 2.895 0.845 3.075 0.855 ;
      RECT 2.895 0.675 3.215 0.845 ;
      RECT 3.045 0.085 3.215 0.675 ;
      RECT 0.785 0.085 1.115 0.94 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 1.805 2.29 2.095 3.245 ;
      RECT 0.645 1.95 1.105 3.245 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a311o_1

MACRO scs8ls_a311o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.55 0.995 2.06 ;
        RECT 0.73 0.75 0.995 1.55 ;
        RECT 0.73 0.35 1.06 0.75 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505 1.45 2.835 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965 1.45 2.295 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.26 1.795 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.26 3.715 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885 1.44 4.215 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END C1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.635 2.57 1.965 2.98 ;
      RECT 1.635 2.29 3.165 2.57 ;
      RECT 2.835 2.57 3.165 2.98 ;
      RECT 1.165 1.95 4.035 2.12 ;
      RECT 3.705 2.12 4.035 2.98 ;
      RECT 1.165 0.92 4.04 1.09 ;
      RECT 3.71 0.35 4.04 0.92 ;
      RECT 2.63 0.35 3 0.92 ;
      RECT 0.105 2.23 1.335 2.4 ;
      RECT 1.165 2.12 1.335 2.23 ;
      RECT 1.165 1.09 1.335 1.95 ;
      RECT 0.105 1.35 0.435 2.23 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 1.23 0.085 1.63 0.75 ;
      RECT 3.17 0.085 3.54 0.75 ;
      RECT 0.3 0.085 0.55 1.13 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 2.135 2.74 2.665 3.245 ;
      RECT 0.215 2.57 0.545 3.245 ;
      RECT 1.115 2.57 1.445 3.245 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a311o_2

MACRO scs8ls_a311o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.45 7.075 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.245 1.45 7.575 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.42 5.295 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535 1.47 1.865 1.8 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.495 1.47 0.825 1.8 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END C1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
    END
  END vpwr

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.095 0.855 2.785 0.995 ;
        RECT 0.095 0.995 0.385 1.04 ;
        RECT 0.095 0.81 0.385 0.855 ;
        RECT 2.495 0.995 2.785 1.04 ;
        RECT 2.495 0.81 2.785 0.855 ;
    END
    ANTENNADIFFAREA 1.0864 ;
    ANTENNAPARTIALMETALSIDEAREA 1.869 LAYER met1 ;
  END X

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 6.285 0.985 7.535 1.245 ;
      RECT 7.285 0.425 7.535 0.985 ;
      RECT 5.365 0.255 7.535 0.425 ;
      RECT 6.775 0.765 7.105 0.815 ;
      RECT 4.415 0.595 7.105 0.765 ;
      RECT 4.415 0.505 4.745 0.595 ;
      RECT 1.735 2.49 1.905 2.735 ;
      RECT 1.735 2.46 5.27 2.49 ;
      RECT 4.94 2.49 5.27 2.98 ;
      RECT 1.735 2.32 6.09 2.46 ;
      RECT 5.92 2.46 6.09 2.98 ;
      RECT 1.735 2.31 1.905 2.32 ;
      RECT 4.94 2.29 6.09 2.32 ;
      RECT 5.92 2.12 6.09 2.29 ;
      RECT 5.92 1.95 7.02 2.12 ;
      RECT 6.85 2.12 7.02 2.98 ;
      RECT 1.205 2.98 2.435 3.075 ;
      RECT 0.305 2.905 2.435 2.98 ;
      RECT 0.305 2.7 1.535 2.905 ;
      RECT 2.105 2.66 2.435 2.905 ;
      RECT 2.535 0.98 3.745 1.15 ;
      RECT 3.495 0.405 3.745 0.98 ;
      RECT 2.535 0.39 2.92 0.98 ;
      RECT 5.545 0.935 6.105 1.265 ;
      RECT 4.475 1.95 5.715 2.12 ;
      RECT 5.545 1.265 5.715 1.95 ;
      RECT 0.905 1.13 2.325 1.3 ;
      RECT 2.055 1.3 2.325 1.32 ;
      RECT 1.755 0.39 1.935 1.13 ;
      RECT 2.055 1.32 3.905 1.48 ;
      RECT 2.055 1.48 4.645 1.65 ;
      RECT 4.475 1.65 4.645 1.95 ;
      RECT 0.755 2.02 1.165 2.19 ;
      RECT 0.995 1.3 1.165 2.02 ;
      RECT 0.905 0.39 1.085 1.13 ;
      RECT 1.335 1.97 4.305 2.14 ;
      RECT 2.525 2.14 4.305 2.15 ;
      RECT 2.525 1.82 4.305 1.97 ;
      RECT 0.125 2.36 1.505 2.53 ;
      RECT 1.335 2.14 1.505 2.36 ;
      RECT 0.125 1.04 0.295 2.36 ;
      RECT 0.125 0.81 0.355 1.04 ;
      RECT 4.175 1.15 5.175 1.185 ;
      RECT 3.925 0.935 5.175 1.15 ;
      RECT 3.925 0.085 4.175 0.935 ;
      RECT 0 -0.085 7.68 0.085 ;
      RECT 0.395 0.085 0.725 0.64 ;
      RECT 1.255 0.085 1.585 0.96 ;
      RECT 2.115 0.085 2.365 0.96 ;
      RECT 3.1 0.085 3.315 0.81 ;
      RECT 0 3.245 7.68 3.415 ;
      RECT 2.625 2.66 2.955 3.245 ;
      RECT 3.525 2.66 3.855 3.245 ;
      RECT 4.425 2.66 4.755 3.245 ;
      RECT 5.47 2.63 5.72 3.245 ;
      RECT 6.29 2.29 6.65 3.245 ;
      RECT 7.22 1.95 7.55 3.245 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 0.84 0.325 1.01 ;
      RECT 2.555 0.84 2.725 1.01 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
  END
END scs8ls_a311o_4

MACRO scs8ls_a311oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 0.35 2.04 1.01 ;
        RECT 0.665 1.01 3.08 1.18 ;
        RECT 0.665 1.18 0.835 1.95 ;
        RECT 2.75 0.35 3.08 1.01 ;
        RECT 0.665 1.95 3.105 2.12 ;
        RECT 2.775 2.12 3.105 2.98 ;
    END
    ANTENNADIFFAREA 0.7927 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.35 1.875 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.35 1.335 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.495 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.35 3.255 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END C1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.765 2.46 1.095 2.98 ;
      RECT 0.765 2.29 2.175 2.46 ;
      RECT 1.845 2.46 2.175 2.98 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 0.34 0.085 0.67 0.84 ;
      RECT 2.21 0.085 2.58 0.84 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 1.265 2.63 1.675 3.245 ;
      RECT 0.315 2.29 0.565 3.245 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a311oi_1

MACRO scs8ls_a311oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.87 1.55 3.235 1.78 ;
        RECT 2.3 1.35 3.235 1.55 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.22 2.09 1.55 ;
        RECT 1.085 1.18 1.315 1.22 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.47 1.22 0.835 1.55 ;
        RECT 0.605 1.18 0.835 1.22 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.35 4.675 1.78 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.845 1.35 5.175 1.78 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END C1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.685 0.35 5.635 1.01 ;
        RECT 2.555 1.01 5.635 1.18 ;
        RECT 5.405 1.18 5.635 1.95 ;
        RECT 2.555 0.85 3.745 1.01 ;
        RECT 4.85 1.95 5.635 2.12 ;
        RECT 3.495 0.35 3.745 0.85 ;
        RECT 4.85 2.12 5.02 2.735 ;
    END
    ANTENNADIFFAREA 0.9354 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.42 2.905 5.55 3.075 ;
      RECT 5.22 2.29 5.55 2.905 ;
      RECT 3.42 2.29 3.755 2.905 ;
      RECT 4.32 1.95 4.65 2.905 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 0.615 0.085 0.945 0.67 ;
      RECT 3.915 0.085 4.515 0.84 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 2.9 2.29 3.23 3.245 ;
      RECT 1.15 2.06 1.32 3.245 ;
      RECT 2.05 2.06 2.33 3.245 ;
      RECT 0.17 1.82 0.42 3.245 ;
      RECT 2.985 0.6 3.315 0.68 ;
      RECT 1.475 0.35 3.315 0.6 ;
      RECT 0.185 1.01 0.435 1.05 ;
      RECT 0.185 0.84 2.235 1.01 ;
      RECT 1.905 1.01 2.235 1.05 ;
      RECT 1.125 0.77 2.235 0.84 ;
      RECT 0.185 0.35 0.435 0.84 ;
      RECT 1.125 0.33 1.295 0.77 ;
      RECT 2.53 1.95 4.12 2.12 ;
      RECT 3.925 2.12 4.12 2.735 ;
      RECT 2.53 2.12 2.7 2.98 ;
      RECT 2.53 1.89 2.7 1.95 ;
      RECT 0.62 1.72 2.7 1.89 ;
      RECT 0.62 1.89 0.95 2.98 ;
      RECT 1.52 1.89 1.85 2.98 ;
    LAYER mcon ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a311oi_2

MACRO scs8ls_a311oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.635 1.35 6.115 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 3.715 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.35 1.875 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.775 1.18 7.555 1.32 ;
        RECT 6.775 1.32 7.785 1.65 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.065 1.22 9.075 1.55 ;
        RECT 8.285 1.18 9.075 1.22 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END C1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.7 0.35 9.955 0.67 ;
        RECT 8.7 0.67 9.425 0.84 ;
        RECT 6.13 0.84 9.425 0.85 ;
        RECT 4.33 0.85 9.425 1.01 ;
        RECT 6.13 0.35 6.38 0.84 ;
        RECT 7.76 0.35 8.01 0.84 ;
        RECT 9.255 1.01 9.425 1.72 ;
        RECT 4.33 1.01 6.38 1.13 ;
        RECT 7.76 1.01 8.01 1.05 ;
        RECT 4.33 0.77 4.66 0.85 ;
        RECT 8.355 1.72 9.425 1.89 ;
        RECT 8.355 1.89 8.525 2.735 ;
        RECT 9.255 1.89 9.425 2.735 ;
    END
    ANTENNADIFFAREA 1.7006 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.3 0.6 2.56 0.68 ;
      RECT 2.3 0.35 5.95 0.6 ;
      RECT 3.23 0.6 3.42 0.68 ;
      RECT 5.62 0.6 5.95 0.68 ;
      RECT 0.15 1.01 3.92 1.18 ;
      RECT 1.95 0.975 3.92 1.01 ;
      RECT 0.15 0.35 0.4 1.01 ;
      RECT 1.01 0.35 1.26 1.01 ;
      RECT 2.73 0.77 3.06 0.975 ;
      RECT 3.59 0.77 3.92 0.975 ;
      RECT 1.95 0.35 2.12 0.975 ;
      RECT 6.525 2.15 6.755 2.735 ;
      RECT 6.475 2.12 7.655 2.15 ;
      RECT 7.425 2.15 7.655 2.735 ;
      RECT 0.555 1.95 7.655 2.12 ;
      RECT 0.555 2.12 0.805 2.98 ;
      RECT 1.535 2.12 1.705 2.98 ;
      RECT 2.435 2.12 2.605 2.98 ;
      RECT 3.335 2.12 3.505 2.98 ;
      RECT 4.235 2.12 4.405 2.98 ;
      RECT 5.055 2.12 5.305 2.98 ;
      RECT 4.235 1.82 4.405 1.95 ;
      RECT 6.475 1.82 7.655 1.95 ;
      RECT 6.025 2.905 9.955 3.075 ;
      RECT 9.625 1.82 9.955 2.905 ;
      RECT 6.025 2.32 6.355 2.905 ;
      RECT 6.925 2.32 7.255 2.905 ;
      RECT 7.825 1.82 8.155 2.905 ;
      RECT 8.725 2.06 9.055 2.905 ;
      RECT 0 -0.085 10.08 0.085 ;
      RECT 0.58 0.085 0.83 0.84 ;
      RECT 1.44 0.085 1.77 0.84 ;
      RECT 6.55 0.085 7.59 0.67 ;
      RECT 8.19 0.085 8.52 0.67 ;
      RECT 0 3.245 10.08 3.415 ;
      RECT 1.005 2.29 1.335 3.245 ;
      RECT 1.905 2.29 2.235 3.245 ;
      RECT 2.805 2.29 3.135 3.245 ;
      RECT 3.705 2.29 4.035 3.245 ;
      RECT 4.605 2.29 4.855 3.245 ;
      RECT 5.505 2.29 5.835 3.245 ;
      RECT 0.105 1.82 0.355 3.245 ;
    LAYER mcon ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
  END
END scs8ls_a311oi_4

MACRO scs8ls_a2111o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.5 2.775 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END D1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.44 0.84 0.67 ;
        RECT 0.51 0.255 0.84 0.44 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.05 1.5 2.275 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.595 0.49 1.795 0.67 ;
        RECT 1.435 0.255 1.795 0.49 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005 0.49 2.245 0.67 ;
        RECT 2.005 0.255 2.335 0.49 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END C1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.86 0.37 4.195 2.98 ;
    END
    ANTENNADIFFAREA 0.5041 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.53 2.14 2.86 2.98 ;
      RECT 2.53 1.97 3.115 2.14 ;
      RECT 2.945 1.65 3.115 1.97 ;
      RECT 2.945 1.33 3.69 1.65 ;
      RECT 0.385 1.32 3.69 1.33 ;
      RECT 0.385 1.16 3.115 1.32 ;
      RECT 2.845 0.66 3.115 1.16 ;
      RECT 1.715 0.84 2.045 1.16 ;
      RECT 0.385 1.33 0.715 1.34 ;
      RECT 0.385 0.84 0.715 1.16 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 2.505 0.085 2.675 0.66 ;
      RECT 3.435 0.085 3.685 1.15 ;
      RECT 2.415 0.66 2.675 0.99 ;
      RECT 1.095 0.66 1.425 0.99 ;
      RECT 1.095 0.085 1.265 0.66 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 0.89 2.31 1.1 3.245 ;
      RECT 3.41 1.82 3.66 3.245 ;
      RECT 0.36 2.14 0.69 2.98 ;
      RECT 0.36 1.97 1.63 2.14 ;
      RECT 1.3 2.14 1.63 2.98 ;
      RECT 0.36 1.94 0.69 1.97 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a2111o_1

MACRO scs8ls_a2111o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.55 0.86 2.98 ;
        RECT 0.69 0.35 0.86 1.55 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.365 1.35 4.695 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.35 4.195 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985 1.35 3.315 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.35 2.775 2.89 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END C1

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.35 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END D1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 1.04 0.085 1.37 0.84 ;
      RECT 2.21 0.085 2.58 0.84 ;
      RECT 3.18 0.085 3.73 0.84 ;
      RECT 0.18 0.085 0.51 1.13 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 3.675 2.29 4.045 3.245 ;
      RECT 1.055 2.29 1.385 3.245 ;
      RECT 0.155 1.82 0.405 3.245 ;
      RECT 3.135 2.12 3.505 2.98 ;
      RECT 3.135 1.95 4.545 2.12 ;
      RECT 4.215 2.12 4.545 2.98 ;
      RECT 1.19 1.01 4.52 1.18 ;
      RECT 4.19 0.35 4.52 1.01 ;
      RECT 2.76 0.35 3.01 1.01 ;
      RECT 1.755 2.12 2.085 2.98 ;
      RECT 1.19 1.95 2.085 2.12 ;
      RECT 1.78 0.35 2.03 1.01 ;
      RECT 1.19 1.55 1.36 1.95 ;
      RECT 1.03 1.22 1.36 1.55 ;
      RECT 1.19 1.18 1.36 1.22 ;
    LAYER mcon ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a2111o_2

MACRO scs8ls_a2111o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.285 1.45 7.075 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.245 1.26 8.035 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405 1.45 6.115 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.45 5.155 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END C1

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385 1.26 3.715 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END D1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.13 0.65 1.8 ;
        RECT 0.125 1.8 2.065 1.97 ;
        RECT 0.125 0.96 2.445 1.13 ;
        RECT 0.835 1.97 1.165 2.98 ;
        RECT 1.735 1.97 2.065 2.98 ;
        RECT 1.415 0.35 1.665 0.96 ;
        RECT 2.195 0.35 2.445 0.96 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 6.01 0.455 6.34 0.94 ;
      RECT 6.01 0.285 7.12 0.455 ;
      RECT 6.95 0.455 7.12 0.92 ;
      RECT 6.95 0.92 8.06 1.09 ;
      RECT 7.81 0.35 8.06 0.92 ;
      RECT 5.025 2.905 6.175 3.075 ;
      RECT 5.025 2.29 5.305 2.905 ;
      RECT 6.005 2.12 6.175 2.905 ;
      RECT 6.005 1.95 8.055 2.12 ;
      RECT 6.905 2.12 7.075 2.98 ;
      RECT 7.725 2.12 8.055 2.98 ;
      RECT 4.135 2.12 4.305 2.735 ;
      RECT 4.135 1.95 5.805 2.12 ;
      RECT 5.475 2.12 5.805 2.735 ;
      RECT 2.705 2.905 4.835 3.075 ;
      RECT 2.705 2.29 3.035 2.905 ;
      RECT 4.505 2.29 4.835 2.905 ;
      RECT 3.605 1.95 3.935 2.905 ;
      RECT 4.05 1.11 6.77 1.28 ;
      RECT 6.51 0.625 6.77 1.11 ;
      RECT 3.045 0.92 4.22 1.09 ;
      RECT 4.05 1.09 4.22 1.11 ;
      RECT 4.05 0.35 4.22 0.92 ;
      RECT 4.92 0.35 5.09 1.11 ;
      RECT 3.235 2.12 3.405 2.735 ;
      RECT 3.045 1.95 3.405 2.12 ;
      RECT 3.045 1.63 3.215 1.95 ;
      RECT 0.87 1.3 3.215 1.63 ;
      RECT 3.045 1.09 3.215 1.3 ;
      RECT 3.045 0.35 3.35 0.92 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 2.625 0.085 2.875 1.03 ;
      RECT 3.53 0.085 3.87 0.75 ;
      RECT 4.4 0.085 4.74 0.94 ;
      RECT 5.27 0.085 5.6 0.94 ;
      RECT 7.3 0.085 7.63 0.75 ;
      RECT 0.905 0.085 1.235 0.79 ;
      RECT 1.845 0.085 2.015 0.79 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 6.375 2.29 6.705 3.245 ;
      RECT 7.275 2.29 7.525 3.245 ;
      RECT 2.265 1.82 2.515 3.245 ;
      RECT 0.385 2.14 0.635 3.245 ;
      RECT 1.365 2.14 1.535 3.245 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
  END
END scs8ls_a2111o_4

MACRO scs8ls_a2111oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.95 1.315 2.98 ;
        RECT 0.125 1.18 0.295 1.95 ;
        RECT 0.125 1.01 2.18 1.18 ;
        RECT 0.85 0.35 1.1 1.01 ;
        RECT 1.85 0.35 2.18 1.01 ;
    END
    ANTENNADIFFAREA 0.7224 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 2.415 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.625 1.18 3.235 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.35 1.875 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.35 1.335 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END C1

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.465 1.35 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END D1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.695 2.12 2.065 2.98 ;
      RECT 1.695 1.95 3.105 2.12 ;
      RECT 2.775 2.12 3.105 2.98 ;
      RECT 2.775 1.82 3.105 1.95 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.75 0.085 3.08 1.01 ;
      RECT 0.34 0.085 0.67 0.84 ;
      RECT 1.27 0.085 1.68 0.84 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.235 2.29 2.605 3.245 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a2111oi_1

MACRO scs8ls_a2111oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.35 4.675 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.85 1.35 5.18 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.35 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END C1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.355 1.95 ;
        RECT 0.125 1.95 1.085 2.12 ;
        RECT 0.125 1.01 2.5 1.18 ;
        RECT 0.755 2.12 1.085 2.735 ;
        RECT 2.17 0.975 2.5 1.01 ;
        RECT 1.16 0.35 1.49 1.01 ;
        RECT 2.17 0.77 4.33 0.975 ;
        RECT 4 0.975 4.33 1.13 ;
        RECT 2.17 0.35 2.5 0.77 ;
    END
    ANTENNADIFFAREA 1.0279 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.18 3.715 1.55 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END B1

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.35 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END D1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.305 2.905 2.435 3.075 ;
      RECT 2.185 2.29 2.435 2.905 ;
      RECT 1.285 1.95 1.455 2.905 ;
      RECT 0.305 2.29 0.555 2.905 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 4.86 0.085 5.2 0.84 ;
      RECT 0.66 0.085 0.99 0.84 ;
      RECT 1.66 0.085 2 0.84 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 4.055 2.29 4.225 3.245 ;
      RECT 4.875 2.29 5.205 3.245 ;
      RECT 4.51 1.01 5.63 1.18 ;
      RECT 4.51 0.6 4.68 1.01 ;
      RECT 5.38 0.35 5.63 1.01 ;
      RECT 3.57 0.35 4.68 0.6 ;
      RECT 2.625 2.905 3.855 3.075 ;
      RECT 2.625 2.29 2.905 2.905 ;
      RECT 3.525 2.12 3.855 2.905 ;
      RECT 3.525 1.95 5.655 2.12 ;
      RECT 4.425 2.12 4.675 2.98 ;
      RECT 5.405 2.12 5.655 2.98 ;
      RECT 5.405 1.82 5.655 1.95 ;
      RECT 1.655 2.12 1.985 2.735 ;
      RECT 1.655 1.95 3.325 2.12 ;
      RECT 3.075 2.12 3.325 2.735 ;
      RECT 3.075 1.82 3.325 1.95 ;
    LAYER mcon ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a2111oi_2

MACRO scs8ls_a2111oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.45 1.35 8.035 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.205 1.35 9.555 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.275 1.35 6.075 1.78 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.235 1.35 3.51 1.78 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END C1

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555 1.18 1.905 1.55 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END D1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.01 0.355 1.72 ;
        RECT 0.125 1.72 1.705 1.89 ;
        RECT 0.125 0.84 2.64 1.01 ;
        RECT 0.555 1.89 0.885 2.735 ;
        RECT 1.455 1.89 1.705 2.735 ;
        RECT 2.39 1.01 7.74 1.13 ;
        RECT 2.39 0.35 2.64 0.84 ;
        RECT 1.53 0.33 1.7 0.84 ;
        RECT 2.39 1.13 6.88 1.18 ;
        RECT 4.07 0.975 7.74 1.01 ;
        RECT 6.55 0.915 7.74 0.975 ;
        RECT 4.07 0.35 4.32 0.975 ;
        RECT 6.55 0.77 6.88 0.915 ;
        RECT 7.41 0.77 7.74 0.915 ;
    END
    ANTENNADIFFAREA 1.708 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 7.92 1.01 9.89 1.18 ;
      RECT 7.92 0.6 8.09 1.01 ;
      RECT 8.78 0.35 8.95 1.01 ;
      RECT 9.64 0.35 9.89 1.01 ;
      RECT 6.12 0.35 8.09 0.6 ;
      RECT 6.12 0.6 6.38 0.68 ;
      RECT 7.04 0.6 7.25 0.68 ;
      RECT 4.245 2.12 4.525 2.735 ;
      RECT 4.245 1.95 9.975 2.12 ;
      RECT 5.195 2.12 5.425 2.735 ;
      RECT 6.125 2.12 6.295 2.98 ;
      RECT 7.025 2.12 7.195 2.98 ;
      RECT 7.925 2.12 8.095 2.98 ;
      RECT 8.745 2.12 9.075 2.98 ;
      RECT 9.725 2.12 9.975 2.98 ;
      RECT 9.725 1.82 9.975 1.95 ;
      RECT 2.435 2.905 5.925 3.075 ;
      RECT 2.435 2.29 2.685 2.905 ;
      RECT 3.255 2.29 3.585 2.905 ;
      RECT 4.695 2.29 5.025 2.905 ;
      RECT 5.595 2.29 5.925 2.905 ;
      RECT 0.105 2.905 2.235 3.075 ;
      RECT 1.905 2.12 2.235 2.905 ;
      RECT 1.905 1.95 4.035 2.12 ;
      RECT 2.855 2.12 3.085 2.735 ;
      RECT 3.755 2.12 4.035 2.735 ;
      RECT 3.705 1.82 4.035 1.95 ;
      RECT 0.105 2.06 0.355 2.905 ;
      RECT 1.085 2.06 1.255 2.905 ;
      RECT 0 -0.085 10.08 0.085 ;
      RECT 8.27 0.085 8.6 0.84 ;
      RECT 9.13 0.085 9.46 0.84 ;
      RECT 1.02 0.085 1.35 0.67 ;
      RECT 1.88 0.085 2.21 0.67 ;
      RECT 2.81 0.085 3.9 0.84 ;
      RECT 4.5 0.085 4.83 0.805 ;
      RECT 0 3.245 10.08 3.415 ;
      RECT 6.495 2.29 6.825 3.245 ;
      RECT 7.395 2.29 7.725 3.245 ;
      RECT 8.295 2.29 8.545 3.245 ;
      RECT 9.275 2.29 9.525 3.245 ;
    LAYER mcon ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
  END
END scs8ls_a2111oi_4

MACRO scs8ls_a211o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.45 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585 1.45 1.835 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 0.255 2.875 0.57 ;
        RECT 2.045 0.57 2.275 0.67 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385 0.255 3.715 0.67 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END C1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.82 0.435 2.98 ;
        RECT 0.085 1.13 0.255 1.82 ;
        RECT 0.085 0.435 1.075 1.13 ;
        RECT 0.825 0.345 1.075 0.435 ;
    END
    ANTENNADIFFAREA 0.5041 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.355 2.12 1.685 2.98 ;
      RECT 1.355 1.95 2.615 2.12 ;
      RECT 2.285 2.12 2.615 2.98 ;
      RECT 1.245 1.11 3.54 1.28 ;
      RECT 3.125 1.28 3.54 2.98 ;
      RECT 2.28 1.08 3.54 1.11 ;
      RECT 2.28 0.84 2.61 1.08 ;
      RECT 0.425 1.4 1.415 1.65 ;
      RECT 1.245 1.28 1.415 1.4 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 2.78 0.74 3.215 0.91 ;
      RECT 3.045 0.085 3.215 0.74 ;
      RECT 1.255 0.085 1.705 0.94 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 1.885 2.29 2.085 3.245 ;
      RECT 0.635 1.82 0.885 3.245 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a211o_1

MACRO scs8ls_a211o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575 1.18 0.835 2.98 ;
        RECT 0.575 1.01 0.98 1.18 ;
        RECT 0.81 0.35 0.98 1.01 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.26 2.535 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.26 1.875 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.745 1.26 3.235 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.45 3.735 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END C1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.545 2.46 1.875 2.98 ;
      RECT 1.545 2.29 2.865 2.46 ;
      RECT 2.535 2.46 2.865 2.98 ;
      RECT 3.405 2.12 3.735 2.98 ;
      RECT 1.165 1.95 3.735 2.12 ;
      RECT 1.165 0.92 3.74 1.09 ;
      RECT 3.49 1.09 3.74 1.13 ;
      RECT 3.49 0.35 3.74 0.92 ;
      RECT 2.33 0.35 2.7 0.92 ;
      RECT 1.165 1.68 1.335 1.95 ;
      RECT 1.005 1.35 1.335 1.68 ;
      RECT 1.165 1.09 1.335 1.35 ;
      RECT 1.16 0.35 1.87 0.75 ;
      RECT 1.16 0.085 1.33 0.35 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 2.87 0.085 3.04 0.35 ;
      RECT 2.87 0.35 3.31 0.75 ;
      RECT 0.3 0.085 0.63 0.84 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 2.075 2.63 2.365 3.245 ;
      RECT 1.025 2.29 1.355 3.245 ;
      RECT 0.125 1.82 0.375 3.245 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a211o_2

MACRO scs8ls_a211o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.45 6.115 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 0.505 5.125 0.67 ;
        RECT 4.925 0.255 5.32 0.505 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.47 4.515 1.72 ;
        RECT 2.785 1.72 4.515 1.89 ;
        RECT 3.995 1.89 4.195 2.15 ;
        RECT 2.785 1.47 3.105 1.72 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.45 1.21 3.78 1.55 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END C1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.33 0.79 2.37 0.96 ;
        RECT 1.33 0.96 1.795 1.24 ;
        RECT 2.18 0.545 2.37 0.79 ;
        RECT 1.33 0.35 1.5 0.79 ;
        RECT 0.675 1.24 1.795 1.41 ;
        RECT 0.675 1.41 0.925 1.72 ;
        RECT 0.675 1.72 1.905 1.89 ;
        RECT 0.675 1.89 0.925 2.98 ;
        RECT 1.575 1.89 1.905 2.98 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 6.235 0.845 6.405 1.275 ;
      RECT 5.295 0.675 6.405 0.845 ;
      RECT 6.235 0.595 6.405 0.675 ;
      RECT 2.545 2.4 4.71 2.57 ;
      RECT 4.5 2.57 4.71 2.99 ;
      RECT 4.42 2.23 4.71 2.4 ;
      RECT 4.42 2.12 5.96 2.23 ;
      RECT 5.725 2.23 5.96 2.98 ;
      RECT 4.42 2.06 6.91 2.12 ;
      RECT 6.63 2.12 6.91 2.98 ;
      RECT 5.68 1.95 6.91 2.06 ;
      RECT 6.58 1.94 6.91 1.95 ;
      RECT 2.545 2.57 2.875 2.78 ;
      RECT 3.96 1.11 6.055 1.28 ;
      RECT 5.725 1.015 6.055 1.11 ;
      RECT 3.04 0.87 4.245 1.04 ;
      RECT 3.96 1.04 4.245 1.11 ;
      RECT 3.96 0.595 4.245 0.87 ;
      RECT 2.445 2.06 3.825 2.23 ;
      RECT 2.445 1.55 2.615 2.06 ;
      RECT 1.965 1.3 2.615 1.55 ;
      RECT 1.965 1.13 3.28 1.3 ;
      RECT 3.04 1.04 3.28 1.13 ;
      RECT 3.04 0.45 3.28 0.87 ;
      RECT 3.045 2.74 4.3 2.99 ;
      RECT 0 -0.085 7.2 0.085 ;
      RECT 6.585 0.085 6.915 1.275 ;
      RECT 3.46 0.085 3.79 0.7 ;
      RECT 4.425 0.085 4.755 0.94 ;
      RECT 2.54 0.085 2.87 0.96 ;
      RECT 0.82 0.085 1.15 1.05 ;
      RECT 1.68 0.085 2.01 0.62 ;
      RECT 0 3.245 7.2 3.415 ;
      RECT 4.88 2.4 5.555 3.245 ;
      RECT 6.13 2.29 6.46 3.245 ;
      RECT 2.105 1.82 2.275 3.245 ;
      RECT 0.225 1.82 0.475 3.245 ;
      RECT 1.125 2.06 1.375 3.245 ;
    LAYER mcon ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
  END
END scs8ls_a211o_4

MACRO scs8ls_a211oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.35 1.335 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.465 1.35 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545 1.35 1.875 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 0.81 2.54 1.01 ;
        RECT 1.085 1.01 2.275 1.025 ;
        RECT 1.085 0.35 1.5 0.81 ;
        RECT 2.21 0.35 2.54 0.81 ;
        RECT 1.085 1.025 2.215 1.18 ;
        RECT 2.045 1.18 2.215 1.82 ;
        RECT 2.045 1.82 2.565 2.98 ;
    END
    ANTENNADIFFAREA 0.7927 ;
  END Y

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.18 2.775 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END C1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.315 2.12 0.645 2.98 ;
      RECT 0.315 1.95 1.635 2.12 ;
      RECT 1.305 2.12 1.635 2.98 ;
      RECT 0 -0.085 2.88 0.085 ;
      RECT 0.34 0.085 0.67 1.13 ;
      RECT 1.67 0.085 2.04 0.64 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 0.815 2.29 1.135 3.245 ;
    LAYER mcon ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a211oi_1

MACRO scs8ls_a211oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.48 1.55 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.43 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.18 3.715 1.55 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.18 4.675 1.55 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END C1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.26 2.755 1.72 ;
        RECT 2.525 1.72 4.145 1.89 ;
        RECT 0.65 1.09 2.755 1.26 ;
        RECT 3.815 1.89 4.145 2.735 ;
        RECT 2.585 1.01 2.755 1.09 ;
        RECT 0.65 0.635 0.83 1.09 ;
        RECT 2.585 0.84 3.59 1.01 ;
        RECT 2.96 0.33 3.59 0.84 ;
    END
    ANTENNADIFFAREA 1.076 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.15 0.255 1.26 0.425 ;
      RECT 1.01 0.425 1.26 0.75 ;
      RECT 1.01 0.75 2.24 0.92 ;
      RECT 1.99 0.33 2.24 0.75 ;
      RECT 0.15 0.425 0.48 1.01 ;
      RECT 1.535 2.12 3.245 2.23 ;
      RECT 2.965 2.23 3.245 2.735 ;
      RECT 0.555 2.06 3.245 2.12 ;
      RECT 1.535 2.23 1.705 2.98 ;
      RECT 0.555 2.12 0.805 2.98 ;
      RECT 0.555 1.95 2.355 2.06 ;
      RECT 0.555 1.82 0.805 1.95 ;
      RECT 2.465 2.905 4.595 3.075 ;
      RECT 4.345 1.82 4.595 2.905 ;
      RECT 2.465 2.4 2.795 2.905 ;
      RECT 3.445 2.06 3.615 2.905 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 3.76 0.085 4.09 1.01 ;
      RECT 1.44 0.33 1.81 0.58 ;
      RECT 1.44 0.085 1.61 0.33 ;
      RECT 2.46 0.085 2.79 0.67 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 1.905 2.4 2.235 3.245 ;
      RECT 1.005 2.29 1.335 3.245 ;
      RECT 0.105 1.82 0.355 3.245 ;
    LAYER mcon ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a211oi_2

MACRO scs8ls_a211oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505 1.35 3.855 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 2.275 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.3 6.115 1.78 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.35 7.555 1.78 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END C1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.18 0.35 8.515 1.01 ;
        RECT 2.57 1.01 8.515 1.13 ;
        RECT 6.32 1.13 8.515 1.18 ;
        RECT 2.57 0.96 6.49 1.01 ;
        RECT 7.725 1.18 8.515 1.95 ;
        RECT 2.57 0.785 3.76 0.96 ;
        RECT 5.38 0.35 5.63 0.96 ;
        RECT 6.32 0.35 6.49 0.96 ;
        RECT 6.795 1.95 7.895 2.12 ;
        RECT 6.795 2.12 6.965 2.735 ;
        RECT 7.695 2.12 7.895 2.735 ;
    END
    ANTENNADIFFAREA 1.6858 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.345 2.12 0.675 2.98 ;
      RECT 0.345 1.95 6.145 2.12 ;
      RECT 1.245 2.12 1.495 2.98 ;
      RECT 2.225 2.12 2.395 2.98 ;
      RECT 3.125 2.12 3.295 2.98 ;
      RECT 4.025 2.12 4.275 2.98 ;
      RECT 4.995 2.12 5.165 2.735 ;
      RECT 5.895 2.12 6.145 2.735 ;
      RECT 4.025 1.82 4.275 1.95 ;
      RECT 2.22 0.35 4.19 0.615 ;
      RECT 0.42 1.01 2.39 1.18 ;
      RECT 2.22 0.615 2.39 1.01 ;
      RECT 0.42 0.35 0.67 1.01 ;
      RECT 1.36 0.35 1.53 1.01 ;
      RECT 4.465 2.905 8.395 3.075 ;
      RECT 8.065 2.12 8.395 2.905 ;
      RECT 4.465 2.29 4.795 2.905 ;
      RECT 5.365 2.29 5.695 2.905 ;
      RECT 6.315 1.95 6.595 2.905 ;
      RECT 7.165 2.29 7.495 2.905 ;
      RECT 0 -0.085 8.64 0.085 ;
      RECT 0.85 0.085 1.18 0.84 ;
      RECT 1.71 0.085 2.04 0.84 ;
      RECT 5.81 0.085 6.14 0.79 ;
      RECT 6.67 0.085 7 0.84 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 0.875 2.29 1.045 3.245 ;
      RECT 1.695 2.29 2.025 3.245 ;
      RECT 2.595 2.29 2.925 3.245 ;
      RECT 3.495 2.29 3.825 3.245 ;
    LAYER mcon ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
  END
END scs8ls_a211oi_4

MACRO scs8ls_a21bo_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.255 0.435 0.67 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.655 1.45 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.515 1.18 2.845 1.55 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END B1N

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.43 1.82 3.755 2.98 ;
        RECT 3.585 1.13 3.755 1.82 ;
        RECT 3.295 0.35 3.755 1.13 ;
    END
    ANTENNADIFFAREA 0.5041 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.13 2.12 0.46 2.98 ;
      RECT 0.13 1.95 1.39 2.12 ;
      RECT 1.06 2.12 1.39 2.98 ;
      RECT 0.13 1.94 0.46 1.95 ;
      RECT 3.085 1.32 3.415 1.65 ;
      RECT 1.575 2.24 3.255 2.41 ;
      RECT 3.085 1.65 3.255 2.24 ;
      RECT 1.575 2.41 1.76 2.98 ;
      RECT 1.575 1.94 1.76 2.24 ;
      RECT 1.575 1.28 1.745 1.94 ;
      RECT 0.945 1.11 1.745 1.28 ;
      RECT 0.945 0.66 1.315 1.11 ;
      RECT 2.075 1.82 2.695 2.07 ;
      RECT 2.075 0.35 2.72 0.94 ;
      RECT 2.075 1.77 2.245 1.82 ;
      RECT 1.915 1.1 2.245 1.77 ;
      RECT 2.075 0.94 2.245 1.1 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 2.9 0.085 3.115 0.895 ;
      RECT 0.155 1.095 0.485 1.34 ;
      RECT 0.155 0.84 0.775 1.095 ;
      RECT 0.605 0.085 0.775 0.84 ;
      RECT 1.485 0.085 1.815 0.93 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 2.9 2.58 3.23 3.245 ;
      RECT 0.66 2.29 0.86 3.245 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a21bo_1

MACRO scs8ls_a21bo_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.02 0.84 1.395 1.04 ;
        RECT 1.225 0.75 1.395 0.84 ;
        RECT 1.02 1.04 1.19 1.82 ;
        RECT 1.225 0.35 1.565 0.75 ;
        RECT 1.02 1.82 1.415 2.07 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.725 1.26 3.235 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.45 3.735 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.51 1.55 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END B1N

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.585 2.27 2.755 2.98 ;
      RECT 2.585 2.1 3.735 2.27 ;
      RECT 3.405 2.27 3.735 2.98 ;
      RECT 3.405 1.95 3.735 2.1 ;
      RECT 1.565 0.92 2.81 1.09 ;
      RECT 2.48 0.35 2.81 0.92 ;
      RECT 2.055 2.06 2.415 2.98 ;
      RECT 2.245 1.93 2.415 2.06 ;
      RECT 2.245 1.76 2.555 1.93 ;
      RECT 2.385 1.09 2.555 1.76 ;
      RECT 1.565 1.09 1.735 1.22 ;
      RECT 1.36 1.22 1.735 1.55 ;
      RECT 0.12 2.24 1.81 2.41 ;
      RECT 1.605 1.89 1.81 2.24 ;
      RECT 1.605 1.72 2.075 1.89 ;
      RECT 1.905 1.59 2.075 1.72 ;
      RECT 1.905 1.26 2.215 1.59 ;
      RECT 0.12 2.41 0.45 2.7 ;
      RECT 0.12 1.82 0.45 2.24 ;
      RECT 0.68 1.01 0.85 2.24 ;
      RECT 0.27 0.84 0.85 1.01 ;
      RECT 0.27 0.54 0.6 0.84 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 1.735 0.085 2.31 0.75 ;
      RECT 3.38 0.085 3.71 1.09 ;
      RECT 0.805 0.085 1.055 0.67 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 0.635 2.58 0.965 3.245 ;
      RECT 1.535 2.58 1.865 3.245 ;
      RECT 2.955 2.44 3.205 3.245 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a21bo_2

MACRO scs8ls_a21bo_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.51 1.42 1.85 ;
        RECT 0.605 1.85 2.3 2.1 ;
        RECT 1.25 1.18 1.42 1.51 ;
        RECT 1.25 1.01 2.415 1.18 ;
        RECT 1.25 0.48 1.555 1.01 ;
        RECT 2.165 0.48 2.415 1.01 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END X

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.45 5.2 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.935 0.255 4.265 0.67 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.505 0.355 0.67 ;
        RECT 0.125 0.255 0.625 0.505 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1N

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.105 2.27 2.64 2.44 ;
      RECT 2.47 2.02 2.64 2.27 ;
      RECT 2.47 1.85 3.29 2.02 ;
      RECT 2.96 1.45 3.29 1.85 ;
      RECT 0.105 2.44 0.435 2.98 ;
      RECT 0.105 1.275 0.435 2.27 ;
      RECT 0.105 0.84 0.615 1.275 ;
      RECT 0 -0.085 6.24 0.085 ;
      RECT 5.725 0.085 5.975 1.275 ;
      RECT 2.595 0.085 2.845 0.94 ;
      RECT 3.595 0.085 3.765 0.94 ;
      RECT 0.795 0.085 1.045 1.275 ;
      RECT 1.735 0.085 1.985 0.84 ;
      RECT 0 3.245 6.24 3.415 ;
      RECT 0.62 2.61 0.95 3.245 ;
      RECT 1.52 2.61 1.85 3.245 ;
      RECT 2.42 2.61 2.75 3.245 ;
      RECT 4.29 2.29 4.54 3.245 ;
      RECT 5.27 2.29 5.52 3.245 ;
      RECT 4.435 0.425 4.605 0.94 ;
      RECT 4.435 0.255 5.545 0.425 ;
      RECT 5.215 0.425 5.545 1.275 ;
      RECT 2.94 2.905 4.09 3.075 ;
      RECT 2.94 2.19 3.27 2.905 ;
      RECT 3.92 2.12 4.09 2.905 ;
      RECT 3.92 1.95 5.97 2.12 ;
      RECT 4.74 2.12 5.07 2.98 ;
      RECT 5.72 2.12 5.97 2.98 ;
      RECT 3.92 1.94 4.09 1.95 ;
      RECT 5.72 1.94 5.97 1.95 ;
      RECT 2.585 1.11 5.035 1.28 ;
      RECT 4.785 0.595 5.035 1.11 ;
      RECT 1.59 1.35 2.755 1.68 ;
      RECT 2.585 1.28 2.755 1.35 ;
      RECT 3.47 1.28 3.72 2.735 ;
      RECT 3.085 0.595 3.415 1.11 ;
    LAYER mcon ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a21bo_4

MACRO scs8ls_a21boi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 2.295 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505 1.18 3.235 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.92 1.525 2.98 ;
        RECT 1.275 1.89 1.525 1.92 ;
        RECT 1.275 1.72 1.875 1.89 ;
        RECT 1.705 1.18 1.875 1.72 ;
        RECT 1.705 1.01 2.06 1.18 ;
        RECT 1.81 0.35 2.06 1.01 ;
    END
    ANTENNADIFFAREA 0.5152 ;
  END Y

  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.12 0.255 0.45 1.605 ;
    END
    ANTENNAGATEAREA 0.208 ;
  END B1N

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.63 0.085 2.96 1.01 ;
      RECT 1.12 0.76 1.45 1.05 ;
      RECT 1.12 0.085 1.63 0.76 ;
      RECT 1.725 2.23 2.02 2.98 ;
      RECT 1.725 2.06 2.985 2.23 ;
      RECT 2.69 2.23 2.985 2.98 ;
      RECT 2.655 1.82 2.985 2.06 ;
      RECT 0.745 1.22 1.535 1.55 ;
      RECT 0.105 1.945 0.435 2.98 ;
      RECT 0.105 1.775 0.915 1.945 ;
      RECT 0.745 1.55 0.915 1.775 ;
      RECT 0.745 1.05 0.95 1.22 ;
      RECT 0.62 0.54 0.95 1.05 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.19 2.4 2.52 3.245 ;
      RECT 0.635 2.115 0.885 3.245 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a21boi_1

MACRO scs8ls_a21boi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.485 1.32 2.815 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.265 1.22 3.715 1.55 ;
        RECT 3.485 1.18 3.715 1.22 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.615 1.15 2.275 1.41 ;
        RECT 1.615 1.41 1.945 2.735 ;
        RECT 1.27 0.98 2.9 1.15 ;
        RECT 2.57 0.77 2.9 0.98 ;
        RECT 1.27 0.35 1.44 0.98 ;
    END
    ANTENNADIFFAREA 0.7504 ;
  END Y

  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.45 0.475 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1N

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.08 1.01 3.25 1.05 ;
      RECT 3.08 0.84 4.19 1.01 ;
      RECT 3.94 1.01 4.19 1.13 ;
      RECT 3.08 0.6 3.25 0.84 ;
      RECT 3.94 0.35 4.19 0.84 ;
      RECT 2.14 0.35 3.25 0.6 ;
      RECT 2.115 1.95 3.215 2.12 ;
      RECT 3.045 2.12 3.215 2.98 ;
      RECT 3.045 1.89 3.215 1.95 ;
      RECT 3.045 1.72 4.215 1.89 ;
      RECT 3.965 1.89 4.215 2.98 ;
      RECT 1.165 2.905 2.315 3.075 ;
      RECT 2.115 2.12 2.315 2.905 ;
      RECT 2.115 1.82 2.315 1.95 ;
      RECT 1.165 1.82 1.415 2.905 ;
      RECT 0.805 1.32 1.395 1.65 ;
      RECT 0.645 1.94 0.975 2.98 ;
      RECT 0.805 1.65 0.975 1.94 ;
      RECT 0.805 1.28 0.975 1.32 ;
      RECT 0.27 1.11 0.975 1.28 ;
      RECT 0.27 0.45 0.52 1.11 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 3.43 0.085 3.76 0.67 ;
      RECT 0.76 0.085 1.09 0.94 ;
      RECT 1.62 0.085 1.95 0.81 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 2.515 2.29 2.845 3.245 ;
      RECT 3.415 2.06 3.765 3.245 ;
      RECT 0.195 1.95 0.445 3.245 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a21boi_2

MACRO scs8ls_a21boi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.43 1.795 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.365 1.43 3.715 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.26 4.745 1.78 ;
        RECT 4.165 1.78 4.745 1.82 ;
        RECT 1.48 1.15 4.745 1.26 ;
        RECT 4.165 1.82 5.395 1.99 ;
        RECT 1.48 1.09 5.72 1.15 ;
        RECT 4.165 1.99 4.495 2.735 ;
        RECT 5.065 1.99 5.395 2.735 ;
        RECT 4.575 0.98 5.72 1.09 ;
        RECT 1.48 0.94 1.81 1.09 ;
        RECT 4.61 0.35 4.86 0.98 ;
        RECT 5.47 0.35 5.72 0.98 ;
        RECT 0.7 0.77 1.81 0.94 ;
        RECT 0.7 0.94 0.95 1.13 ;
    END
    ANTENNADIFFAREA 1.5008 ;
  END Y

  PIN B1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.49 7.555 1.82 ;
    END
    ANTENNAGATEAREA 0.363 ;
  END B1N

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.19 0.35 2.16 0.6 ;
      RECT 1.99 0.6 2.16 0.75 ;
      RECT 1.99 0.75 3.96 0.92 ;
      RECT 2.85 0.51 3.02 0.75 ;
      RECT 3.71 0.51 3.96 0.75 ;
      RECT 0.19 0.6 0.52 1.13 ;
      RECT 3.715 2.905 5.845 3.075 ;
      RECT 5.565 1.82 5.845 2.905 ;
      RECT 3.715 2.12 3.995 2.905 ;
      RECT 0.115 1.95 3.995 2.12 ;
      RECT 0.115 2.12 0.365 2.98 ;
      RECT 1.095 2.12 1.265 2.98 ;
      RECT 1.995 2.12 2.165 2.98 ;
      RECT 2.815 2.12 3.145 2.98 ;
      RECT 1.995 1.82 2.165 1.95 ;
      RECT 4.665 2.16 4.895 2.905 ;
      RECT 6.535 2.16 6.815 2.98 ;
      RECT 6.025 1.99 6.815 2.16 ;
      RECT 6.025 1.15 6.66 1.32 ;
      RECT 6.4 0.35 6.66 1.15 ;
      RECT 6.025 1.65 6.195 1.99 ;
      RECT 4.915 1.32 6.195 1.65 ;
      RECT 0 -0.085 7.68 0.085 ;
      RECT 5.9 0.085 6.23 0.98 ;
      RECT 2.34 0.085 2.67 0.58 ;
      RECT 3.2 0.085 3.53 0.58 ;
      RECT 4.18 0.085 4.43 0.88 ;
      RECT 5.04 0.085 5.29 0.81 ;
      RECT 0 3.245 7.68 3.415 ;
      RECT 6.035 2.33 6.365 3.245 ;
      RECT 7.015 2.1 7.265 3.245 ;
      RECT 0.565 2.29 0.895 3.245 ;
      RECT 1.465 2.29 1.795 3.245 ;
      RECT 2.365 2.29 2.615 3.245 ;
      RECT 3.345 2.29 3.515 3.245 ;
    LAYER mcon ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
  END
END scs8ls_a21boi_4

MACRO scs8ls_a21o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.645 0.255 3.235 0.57 ;
        RECT 3.005 0.57 3.235 0.67 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585 1.45 1.835 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.45 2.375 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.82 0.435 2.98 ;
        RECT 0.085 1.15 0.255 1.82 ;
        RECT 0.085 0.98 1.075 1.15 ;
        RECT 0.825 0.67 1.075 0.98 ;
    END
    ANTENNADIFFAREA 0.5041 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.805 2.12 2.135 2.98 ;
      RECT 1.805 1.95 3.065 2.12 ;
      RECT 2.735 2.12 3.065 2.98 ;
      RECT 2.735 1.94 3.065 1.95 ;
      RECT 1.245 1.11 2.135 1.28 ;
      RECT 1.805 0.66 2.135 1.11 ;
      RECT 1.245 1.95 1.605 2.98 ;
      RECT 1.245 1.65 1.415 1.95 ;
      RECT 0.425 1.32 1.415 1.65 ;
      RECT 1.245 1.28 1.415 1.32 ;
      RECT 2.71 1.01 3.04 1.34 ;
      RECT 2.305 0.84 3.04 1.01 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.305 0.085 2.475 0.84 ;
      RECT 1.255 0.085 1.585 0.94 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.335 2.29 2.535 3.245 ;
      RECT 0.635 1.82 0.885 3.245 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a21o_1

MACRO scs8ls_a21o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.57 1.55 0.9 1.89 ;
        RECT 0.57 1.89 0.85 2.98 ;
        RECT 0.725 1.05 0.9 1.55 ;
        RECT 0.725 0.35 1.055 1.05 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.2 1.18 2.755 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.18 3.255 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.18 1.99 1.535 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.99 1.89 2.24 2.98 ;
      RECT 1.99 1.72 3.22 1.89 ;
      RECT 2.97 1.89 3.22 2.98 ;
      RECT 1.225 0.84 2.295 1.01 ;
      RECT 1.965 0.35 2.295 0.84 ;
      RECT 1.54 1.875 1.79 2.98 ;
      RECT 1.07 1.705 1.79 1.875 ;
      RECT 1.07 1.22 1.395 1.705 ;
      RECT 1.225 1.01 1.395 1.22 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 1.225 0.085 1.795 0.67 ;
      RECT 2.865 0.085 3.195 1.01 ;
      RECT 0.295 0.085 0.545 1.13 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.44 2.06 2.77 3.245 ;
      RECT 1.02 2.045 1.35 3.245 ;
      RECT 0.12 1.82 0.37 3.245 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a21o_2

MACRO scs8ls_a21o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.45 4.195 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.26 4.905 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.425 1.435 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.492 ;
  END B1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.13 0.355 1.8 ;
        RECT 0.125 1.8 1.835 1.97 ;
        RECT 0.125 0.96 1.69 1.13 ;
        RECT 0.685 1.97 0.855 2.98 ;
        RECT 1.505 1.97 1.835 2.98 ;
        RECT 0.66 0.35 0.83 0.96 ;
        RECT 1.44 0.35 1.69 0.96 ;
    END
    ANTENNADIFFAREA 1.0864 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 3.825 2.29 4.075 3.245 ;
      RECT 4.725 2.29 5.055 3.245 ;
      RECT 2.035 1.95 2.285 3.245 ;
      RECT 0.155 2.14 0.485 3.245 ;
      RECT 1.055 2.14 1.305 3.245 ;
      RECT 3.46 0.425 3.79 0.94 ;
      RECT 3.46 0.255 4.57 0.425 ;
      RECT 4.4 0.425 4.57 0.92 ;
      RECT 4.4 0.92 5.51 1.09 ;
      RECT 5.26 0.35 5.51 0.92 ;
      RECT 2.475 2.905 3.625 3.075 ;
      RECT 3.455 2.12 3.625 2.905 ;
      RECT 2.475 1.95 2.725 2.905 ;
      RECT 3.455 1.95 5.505 2.12 ;
      RECT 4.275 2.12 4.525 2.98 ;
      RECT 5.255 2.12 5.505 2.98 ;
      RECT 5.255 1.94 5.505 1.95 ;
      RECT 1.87 1.11 4.22 1.265 ;
      RECT 2.925 1.265 4.22 1.28 ;
      RECT 3.96 0.595 4.22 1.11 ;
      RECT 1.87 1.095 3.255 1.11 ;
      RECT 2.925 1.28 3.255 2.735 ;
      RECT 2.36 0.45 2.61 1.095 ;
      RECT 0.635 1.3 2.205 1.63 ;
      RECT 1.87 1.265 2.205 1.3 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 1.87 0.085 2.12 0.925 ;
      RECT 2.79 0.085 3.12 0.925 ;
      RECT 4.75 0.085 5.08 0.75 ;
      RECT 0.15 0.085 0.48 0.79 ;
      RECT 1.01 0.085 1.26 0.79 ;
    LAYER mcon ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a21o_4

MACRO scs8ls_a21oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.35 1.05 1.78 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.18 0.435 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.89 1.815 2.98 ;
        RECT 1.22 1.72 1.815 1.89 ;
        RECT 1.22 1.18 1.39 1.72 ;
        RECT 0.92 1.01 1.39 1.18 ;
        RECT 0.92 0.35 1.29 1.01 ;
    END
    ANTENNADIFFAREA 0.5966 ;
  END Y

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.56 1.19 1.815 1.55 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END B1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.105 2.06 1.365 2.23 ;
      RECT 1.07 2.23 1.365 2.98 ;
      RECT 0.105 2.23 0.4 2.98 ;
      RECT 0.105 1.985 0.955 2.06 ;
      RECT 0.105 1.82 0.435 1.985 ;
      RECT 0 -0.085 1.92 0.085 ;
      RECT 1.56 0.085 1.79 1.02 ;
      RECT 0.13 0.085 0.46 1.01 ;
      RECT 0 3.245 1.92 3.415 ;
      RECT 0.57 2.4 0.9 3.245 ;
    LAYER mcon ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a21oi_1

MACRO scs8ls_a21oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.35 3.35 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.18 2.755 1.78 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.435 0.435 1.78 ;
    END
    ANTENNAGATEAREA 0.447 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.55 1.395 1.78 ;
        RECT 1.065 1.78 1.395 2.735 ;
        RECT 0.605 0.92 0.86 1.55 ;
        RECT 0.605 0.75 3.18 0.92 ;
        RECT 2.93 0.92 3.18 1.13 ;
        RECT 0.605 0.35 0.86 0.75 ;
    END
    ANTENNADIFFAREA 0.7393 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.615 2.905 1.845 3.075 ;
      RECT 1.565 2.46 1.845 2.905 ;
      RECT 1.565 2.29 3.705 2.46 ;
      RECT 2.475 2.46 2.805 2.98 ;
      RECT 3.375 2.46 3.705 2.98 ;
      RECT 0.615 1.95 0.895 2.905 ;
      RECT 1.565 1.95 3.69 2.12 ;
      RECT 3.52 1.13 3.69 1.95 ;
      RECT 3.36 0.58 3.69 1.13 ;
      RECT 2.5 0.33 3.69 0.58 ;
      RECT 1.565 1.26 1.775 1.95 ;
      RECT 1.36 1.09 1.775 1.26 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 0.1 0.085 0.43 1.13 ;
      RECT 2 0.085 2.33 0.58 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 2.045 2.63 2.305 3.245 ;
      RECT 3.005 2.63 3.175 3.245 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a21oi_2

MACRO scs8ls_a21oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 1.35 3.935 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.785 1.35 2.275 1.78 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.235 1.35 5.245 1.78 ;
    END
    ANTENNAGATEAREA 0.894 ;
  END B1

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 0.88 4.65 1.01 ;
        RECT 2.525 1.01 5.59 1.18 ;
        RECT 2.525 0.595 2.78 0.88 ;
        RECT 4.4 0.35 4.65 0.88 ;
        RECT 2.525 1.18 2.755 1.95 ;
        RECT 5.34 0.35 5.59 1.01 ;
        RECT 2.525 1.95 5.585 2.12 ;
        RECT 4.355 2.12 4.685 2.735 ;
        RECT 5.255 2.12 5.585 2.735 ;
    END
    ANTENNADIFFAREA 1.4786 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.905 2.905 6.035 3.075 ;
      RECT 5.785 1.82 6.035 2.905 ;
      RECT 2.105 2.46 2.355 2.98 ;
      RECT 2.105 2.12 2.355 2.29 ;
      RECT 0.305 1.95 2.355 2.12 ;
      RECT 0.305 2.12 0.555 2.98 ;
      RECT 1.205 2.12 1.535 2.98 ;
      RECT 0.305 1.82 0.555 1.95 ;
      RECT 2.105 2.29 4.155 2.46 ;
      RECT 3.005 2.46 3.335 2.98 ;
      RECT 3.905 2.46 4.155 2.905 ;
      RECT 4.885 2.29 5.055 2.905 ;
      RECT 0 -0.085 6.24 0.085 ;
      RECT 0.81 0.085 1.14 0.84 ;
      RECT 1.67 0.085 2 0.84 ;
      RECT 4.83 0.085 5.16 0.84 ;
      RECT 0 3.245 6.24 3.415 ;
      RECT 2.555 2.63 2.805 3.245 ;
      RECT 3.535 2.63 3.705 3.245 ;
      RECT 0.755 2.29 1.005 3.245 ;
      RECT 1.735 2.29 1.905 3.245 ;
      RECT 2.18 0.255 4.15 0.425 ;
      RECT 2.96 0.425 3.29 0.71 ;
      RECT 3.82 0.425 4.15 0.71 ;
      RECT 0.38 1.01 2.35 1.18 ;
      RECT 2.18 0.425 2.35 1.01 ;
      RECT 0.38 0.35 0.63 1.01 ;
      RECT 1.32 0.35 1.49 1.01 ;
    LAYER mcon ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a21oi_4

MACRO scs8ls_a221o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.455 2.985 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B1

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965 1.47 2.295 1.8 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.375 1.35 1.795 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END A2

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.195 1.455 3.715 1.78 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.865 0.255 4.195 0.67 ;
    END
    ANTENNAGATEAREA 0.246 ;
  END C1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.82 0.9 2.98 ;
        RECT 0.125 1.13 0.5 1.82 ;
        RECT 0.125 0.35 0.865 1.13 ;
    END
    ANTENNADIFFAREA 0.5041 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.535 2.14 1.785 2.98 ;
      RECT 1.535 1.97 3.285 2.14 ;
      RECT 2.955 2.14 3.285 2.735 ;
      RECT 1.535 1.95 1.785 1.97 ;
      RECT 2.955 1.95 3.285 1.97 ;
      RECT 2.505 2.905 3.685 3.075 ;
      RECT 2.505 2.31 2.785 2.905 ;
      RECT 3.485 1.95 3.685 2.905 ;
      RECT 1.035 1.115 4.215 1.18 ;
      RECT 2.465 1.18 4.215 1.285 ;
      RECT 3.86 0.84 4.215 1.115 ;
      RECT 3.885 1.285 4.215 2.98 ;
      RECT 1.035 1.01 2.86 1.115 ;
      RECT 2.42 0.375 2.86 1.01 ;
      RECT 0.74 1.3 1.205 1.63 ;
      RECT 1.035 1.18 1.205 1.3 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 1.045 0.085 1.965 0.84 ;
      RECT 3.32 0.085 3.69 0.945 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 1.985 2.31 2.315 3.245 ;
      RECT 1.1 1.95 1.35 3.245 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a221o_1

MACRO scs8ls_a221o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.32 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.6 1.97 0.93 2.98 ;
        RECT 0.1 1.8 0.93 1.97 ;
        RECT 0.1 1.13 0.335 1.8 ;
        RECT 0.1 0.96 0.855 1.13 ;
        RECT 0.605 0.35 0.855 0.96 ;
    END
    ANTENNADIFFAREA 0.5432 ;
  END X

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935 1.45 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.365 1.26 1.765 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.455 1.45 2.76 1.78 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.27 1.18 3.695 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.865 1.18 4.195 1.55 ;
    END
    ANTENNAGATEAREA 0.261 ;
  END C1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.32 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.32 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.985 2.23 3.315 2.735 ;
      RECT 2.54 2.12 3.315 2.23 ;
      RECT 1.565 2.06 3.315 2.12 ;
      RECT 1.565 2.12 1.815 2.98 ;
      RECT 1.565 1.95 2.73 2.06 ;
      RECT 2.535 2.905 3.685 3.075 ;
      RECT 2.535 2.4 2.785 2.905 ;
      RECT 3.515 2.06 3.685 2.905 ;
      RECT 3.885 1.89 4.215 2.98 ;
      RECT 2.93 1.72 4.215 1.89 ;
      RECT 1.025 0.92 4.22 1.01 ;
      RECT 2.02 0.84 4.22 0.92 ;
      RECT 3.89 0.35 4.22 0.84 ;
      RECT 2.93 1.13 3.1 1.72 ;
      RECT 2.02 1.09 3.1 1.13 ;
      RECT 1.025 1.01 3.1 1.09 ;
      RECT 2.02 0.35 2.89 0.84 ;
      RECT 1.025 1.09 1.195 1.3 ;
      RECT 0.525 1.3 1.195 1.63 ;
      RECT 0 -0.085 4.32 0.085 ;
      RECT 1.035 0.085 1.56 0.75 ;
      RECT 3.35 0.085 3.72 0.67 ;
      RECT 0.175 0.085 0.425 0.79 ;
      RECT 0 3.245 4.32 3.415 ;
      RECT 2.015 2.29 2.345 3.245 ;
      RECT 1.13 1.95 1.38 3.245 ;
      RECT 0.15 2.14 0.4 3.245 ;
    LAYER mcon ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_a221o_2


MACRO scs8ls_probe_s8p_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.43 1.78 ;
    END
    ANTENNAGATEAREA 0.837 LAYER met1 ;
    ANTENNAGATEAREA 0.837 LAYER met2 ;
    ANTENNAGATEAREA 0.837 LAYER met3 ;
    ANTENNAGATEAREA 0.837 LAYER met4 ;
    ANTENNAGATEAREA 0.837 LAYER met5 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1.37 0.865 4.39 2.465 ;
    END
    PORT
      LAYER via4 ;
        RECT 1.68 1.175 2.48 1.975 ;
        RECT 3.28 1.175 4.08 1.975 ;
    END
    ANTENNAPARTIALMETALSIDEAREA 0.02 LAYER met5 ;
  END X

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met4 ;
      RECT 1.49 0.985 4.27 2.165 ;
      RECT 3.54 1.4 4.27 1.73 ;
    LAYER met3 ;
      RECT 3.54 1.4 4.27 1.73 ;
      RECT 3.515 1.405 4.295 1.725 ;
      RECT 3.515 1.4 3.54 1.73 ;
      RECT 4.27 1.4 4.295 1.73 ;
    LAYER met2 ;
      RECT 3.585 1.435 4.225 1.695 ;
      RECT 3.565 1.38 4.245 1.75 ;
    LAYER met1 ;
      RECT 3.585 1.435 4.225 1.695 ;
      RECT 4.225 1.45 4.745 1.68 ;
      RECT 4.745 1.45 5.395 1.68 ;
    LAYER li1 ;
      RECT 1.97 1.97 2.3 2.98 ;
      RECT 1.97 1.8 5.155 1.97 ;
      RECT 2.92 1.97 3.25 2.98 ;
      RECT 3.87 1.97 4.2 2.98 ;
      RECT 4.82 1.97 5.155 2.98 ;
      RECT 4.805 1.13 5.145 1.48 ;
      RECT 4.805 1.48 5.335 1.65 ;
      RECT 1.96 0.96 5.145 1.13 ;
      RECT 1.96 0.35 2.13 0.96 ;
      RECT 2.81 0.35 3.14 0.96 ;
      RECT 3.81 0.35 4.14 0.96 ;
      RECT 4.81 0.35 5.145 0.96 ;
      RECT 4.805 1.65 5.155 1.8 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 0.65 2.29 0.82 3.245 ;
      RECT 1.55 2.29 1.8 3.245 ;
      RECT 2.5 2.14 2.75 3.245 ;
      RECT 3.45 2.14 3.7 3.245 ;
      RECT 4.4 2.14 4.65 3.245 ;
      RECT 5.35 1.82 5.6 3.245 ;
      RECT 0.545 0.085 0.875 0.84 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 1.45 0.085 1.78 0.84 ;
      RECT 2.31 0.085 2.64 0.79 ;
      RECT 3.31 0.085 3.64 0.79 ;
      RECT 4.31 0.085 4.64 0.79 ;
      RECT 5.315 0.085 5.645 1.13 ;
      RECT 0.12 2.12 0.45 2.98 ;
      RECT 0.12 1.95 1.77 2.12 ;
      RECT 1.02 2.12 1.35 2.98 ;
      RECT 1.6 1.63 1.77 1.95 ;
      RECT 1.6 1.3 4.605 1.63 ;
      RECT 1.6 1.18 1.77 1.3 ;
      RECT 0.115 1.01 1.77 1.18 ;
      RECT 0.115 0.35 0.365 1.01 ;
      RECT 1.1 0.35 1.27 1.01 ;
    LAYER via3 ;
      RECT 4.005 1.465 4.205 1.665 ;
      RECT 3.605 1.465 3.805 1.665 ;
    LAYER via2 ;
      RECT 3.605 1.465 3.805 1.665 ;
      RECT 4.005 1.465 4.205 1.665 ;
    LAYER via ;
      RECT 3.99 1.49 4.14 1.64 ;
      RECT 3.67 1.49 3.82 1.64 ;
    LAYER mcon ;
      RECT 4.805 1.48 4.975 1.65 ;
      RECT 5.165 1.48 5.335 1.65 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_probe_s8p_8

MACRO scs8ls_probec_s8p_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.43 1.78 ;
    END
    ANTENNAGATEAREA 0.837 LAYER met1 ;
    ANTENNAGATEAREA 0.837 LAYER met2 ;
    ANTENNAGATEAREA 0.837 LAYER met3 ;
    ANTENNAGATEAREA 0.837 LAYER met4 ;
    ANTENNAGATEAREA 0.837 LAYER met5 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.13 6.08 0.13 ;
        RECT 0 0.13 5.76 0.245 ;
        RECT 0 -0.245 5.76 -0.13 ;
    END
    PORT
      LAYER via ;
        RECT 5.845 -0.075 5.995 0.075 ;
        RECT 5.525 -0.075 5.675 0.075 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.2 6.08 3.46 ;
        RECT 0 3.46 5.76 3.575 ;
        RECT 0 3.085 5.76 3.2 ;
    END
    PORT
      LAYER via ;
        RECT 5.525 3.255 5.675 3.405 ;
        RECT 5.845 3.255 5.995 3.405 ;
    END
  END vpwr

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -0.475 1.505 0.305 1.825 ;
    END
    PORT
      LAYER via3 ;
        RECT -0.385 1.565 -0.185 1.765 ;
        RECT 0.015 1.565 0.215 1.765 ;
    END
    ANTENNAPARTIALMETALSIDEAREA 0.736 LAYER met3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.776 LAYER met4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.32 LAYER met5 ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3 ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4 ;
  END X

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met5 ;
      RECT 4.6 2.465 6.915 4.195 ;
      RECT 4.6 -0.865 6.915 0.865 ;
      RECT -1.02 0.865 3 2.465 ;
      RECT 1.4 2.465 3 4.13 ;
      RECT 1.4 -0.8 3 0.865 ;
    LAYER met4 ;
      RECT 5.17 -0.59 6.35 0.59 ;
      RECT 5.17 2.74 6.35 3.92 ;
      RECT 1.7 1.075 2.88 2.255 ;
      RECT -0.9 1.075 0.28 2.255 ;
    LAYER met3 ;
      RECT 5.37 -0.165 6.15 0.165 ;
      RECT 5.37 3.165 6.15 3.495 ;
      RECT 2.125 1.5 2.905 1.83 ;
    LAYER met2 ;
      RECT 5.375 -0.14 6.145 0.14 ;
      RECT 5.375 3.19 6.145 3.47 ;
      RECT 2.13 1.525 2.9 1.805 ;
      RECT 2.26 1.435 2.9 1.525 ;
    LAYER met1 ;
      RECT 2.26 1.435 2.9 1.695 ;
      RECT 2.26 1.45 4.745 1.68 ;
      RECT 4.745 1.45 5.395 1.68 ;
    LAYER li1 ;
      RECT 1.97 1.97 2.3 2.98 ;
      RECT 1.97 1.8 5.155 1.97 ;
      RECT 2.92 1.97 3.25 2.98 ;
      RECT 3.87 1.97 4.2 2.98 ;
      RECT 4.82 1.97 5.155 2.98 ;
      RECT 4.805 1.13 5.145 1.48 ;
      RECT 4.805 1.48 5.335 1.65 ;
      RECT 1.96 0.96 5.145 1.13 ;
      RECT 1.96 0.35 2.13 0.96 ;
      RECT 2.81 0.35 3.14 0.96 ;
      RECT 3.81 0.35 4.14 0.96 ;
      RECT 4.81 0.35 5.145 0.96 ;
      RECT 4.805 1.65 5.155 1.8 ;
      RECT 0.545 0.085 0.875 0.84 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 1.45 0.085 1.78 0.84 ;
      RECT 2.31 0.085 2.64 0.79 ;
      RECT 3.31 0.085 3.64 0.79 ;
      RECT 4.31 0.085 4.64 0.79 ;
      RECT 5.315 0.085 5.645 1.13 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 0.65 2.29 0.82 3.245 ;
      RECT 1.55 2.29 1.8 3.245 ;
      RECT 2.5 2.14 2.75 3.245 ;
      RECT 3.45 2.14 3.7 3.245 ;
      RECT 4.4 2.14 4.65 3.245 ;
      RECT 5.35 1.82 5.6 3.245 ;
      RECT 0.12 2.12 0.45 2.98 ;
      RECT 0.12 1.95 1.77 2.12 ;
      RECT 1.02 2.12 1.35 2.98 ;
      RECT 1.6 1.63 1.77 1.95 ;
      RECT 1.6 1.3 4.605 1.63 ;
      RECT 1.6 1.18 1.77 1.3 ;
      RECT 0.115 1.01 1.77 1.18 ;
      RECT 0.115 0.35 0.365 1.01 ;
      RECT 1.1 0.35 1.27 1.01 ;
    LAYER via4 ;
      RECT 5.36 -0.4 6.16 0.4 ;
      RECT 5.36 2.93 6.16 3.73 ;
      RECT 1.89 1.265 2.69 2.065 ;
      RECT -0.71 1.265 0.09 2.065 ;
    LAYER via3 ;
      RECT 5.86 -0.1 6.06 0.1 ;
      RECT 5.46 -0.1 5.66 0.1 ;
      RECT 5.46 3.23 5.66 3.43 ;
      RECT 5.86 3.23 6.06 3.43 ;
      RECT 2.215 1.565 2.415 1.765 ;
      RECT 2.615 1.565 2.815 1.765 ;
    LAYER via2 ;
      RECT 5.46 -0.1 5.66 0.1 ;
      RECT 5.86 -0.1 6.06 0.1 ;
      RECT 5.46 3.23 5.66 3.43 ;
      RECT 5.86 3.23 6.06 3.43 ;
      RECT 2.215 1.565 2.415 1.765 ;
      RECT 2.615 1.565 2.815 1.765 ;
    LAYER via ;
      RECT 2.345 1.49 2.495 1.64 ;
      RECT 2.665 1.49 2.815 1.64 ;
    LAYER mcon ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 4.805 1.48 4.975 1.65 ;
      RECT 5.165 1.48 5.335 1.65 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
  END
END scs8ls_probec_s8p_8

  
END LIBRARY
