# 
# LEF OUT 
# User Name : apoe 
# Date : Thu Jun  4 08:27:35 2020
# 
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO scs8ls_udb_tapmet1_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.96 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.96 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.56 2.645 0.88 2.905 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.08 0.425 0.4 0.685 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.09 0.265 0.87 1.105 ;
      RECT 0 -0.085 0.96 0.085 ;
      RECT 0 3.245 0.96 3.415 ;
      RECT 0.09 2.21 0.87 3.065 ;
    LAYER mcon ;
      RECT 0.635 2.69 0.805 2.86 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 0.47 0.325 0.64 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_udb_tapmet1_2

MACRO scs8ls_udb_a2222o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.76 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.325 1.165 5.655 1.495 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END A2

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.465 1.165 3.795 1.495 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END B2

  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995 1.165 1.325 1.495 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END D2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.65 1.165 5.155 1.495 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.099 LAYER li1 ;
  END A1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.165 4.44 1.495 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.093 LAYER li1 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.065 1.165 2.595 1.495 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.104 LAYER li1 ;
  END C1

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.82 0.365 2.98 ;
        RECT 0.085 1.13 0.255 1.82 ;
        RECT 0.085 0.35 0.445 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
    ANTENNAPARTIALMETALSIDEAREA 0.416 LAYER li1 ;
  END X

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.165 1.895 1.495 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END D1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.805 1.165 3.235 1.495 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER li1 ;
  END C2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.76 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.76 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.515 2.61 3.845 2.98 ;
      RECT 3.515 2.44 4.665 2.61 ;
      RECT 4.495 2.61 4.665 2.98 ;
      RECT 4.495 1.835 4.665 2.44 ;
      RECT 4.495 1.665 5.645 1.835 ;
      RECT 5.395 1.835 5.645 2.98 ;
      RECT 2.475 1.94 4.295 2.27 ;
      RECT 1.125 2.61 1.455 2.98 ;
      RECT 1.125 2.44 3.285 2.61 ;
      RECT 2.025 2.61 2.355 2.98 ;
      RECT 2.955 2.61 3.285 2.98 ;
      RECT 0.615 0.825 4.485 0.995 ;
      RECT 4.235 0.35 4.485 0.825 ;
      RECT 1.69 0.665 2.44 0.825 ;
      RECT 1.575 1.835 1.905 2.27 ;
      RECT 0.615 1.665 1.905 1.835 ;
      RECT 0.615 1.63 0.785 1.665 ;
      RECT 0.425 1.3 0.785 1.63 ;
      RECT 0.615 0.995 0.785 1.3 ;
      RECT 0.625 0.085 1.12 0.655 ;
      RECT 0 -0.085 5.76 0.085 ;
      RECT 3.01 0.085 3.665 0.655 ;
      RECT 5.395 0.085 5.645 0.995 ;
      RECT 0 3.245 5.76 3.415 ;
      RECT 0.565 2.005 0.895 3.245 ;
      RECT 4.865 2.005 5.195 3.245 ;
    LAYER mcon ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_udb_a2222o_1

MACRO scs8ls_udb_a2222o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.35 4.305 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.086 LAYER li1 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.805 1.3 6.135 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.094 LAYER li1 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.475 1.45 4.895 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.082 LAYER li1 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.105 1.45 5.635 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.104 LAYER li1 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455 1.47 1.795 1.8 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.066 LAYER li1 ;
  END C1

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.99 1.45 1.285 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.057 LAYER li1 ;
  END D1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.995 1.18 2.325 1.8 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.054 LAYER li1 ;
  END C2

  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.45 0.48 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.069 LAYER li1 ;
  END D2

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.45 1.55 3.715 1.82 ;
        RECT 3.335 1.82 3.715 2.07 ;
        RECT 3.45 1.09 3.62 1.55 ;
        RECT 2.835 0.92 3.62 1.09 ;
    END
    ANTENNADIFFAREA 0.6172 ;
    ANTENNAPARTIALMETALSIDEAREA 0.361 LAYER li1 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.79 0.96 6.125 1.13 ;
      RECT 3.79 0.92 4.23 0.96 ;
      RECT 5.875 0.46 6.125 0.96 ;
      RECT 4.29 2.75 4.62 2.98 ;
      RECT 4.29 2.58 5.625 2.75 ;
      RECT 5.295 2.75 5.625 2.98 ;
      RECT 5.295 1.95 5.625 2.58 ;
      RECT 1.645 2.24 5.125 2.41 ;
      RECT 4.79 2.08 5.125 2.24 ;
      RECT 1.645 2.41 1.975 2.735 ;
      RECT 1.645 1.97 1.975 2.24 ;
      RECT 0.145 2.905 2.665 3.075 ;
      RECT 2.145 2.65 2.665 2.905 ;
      RECT 1.145 1.97 1.475 2.905 ;
      RECT 0.145 1.95 0.475 2.905 ;
      RECT 1.04 0.58 4.685 0.75 ;
      RECT 4.33 0.5 4.685 0.58 ;
      RECT 2.495 0.75 2.665 1.26 ;
      RECT 0.65 1.11 1.37 1.28 ;
      RECT 1.04 0.75 1.37 1.11 ;
      RECT 0.645 1.95 0.975 2.735 ;
      RECT 0.65 1.28 0.82 1.95 ;
      RECT 2.495 1.26 3.28 1.59 ;
      RECT 5.26 0.46 5.695 0.79 ;
      RECT 5.525 0.085 5.695 0.46 ;
      RECT 0 -0.085 6.24 0.085 ;
      RECT 3.345 0.085 3.705 0.41 ;
      RECT 2.135 0.085 2.555 0.4 ;
      RECT 0.15 0.085 0.48 1.28 ;
      RECT 0 3.245 6.24 3.415 ;
      RECT 3.785 2.58 4.115 3.245 ;
      RECT 5.795 1.95 6.125 3.245 ;
      RECT 2.885 2.58 3.215 3.245 ;
    LAYER mcon ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_udb_a2222o_2

MACRO scs8ls_udb_a2222oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.845 1.3 5.175 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.094 LAYER li1 ;
  END A2

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.92 1.45 3.25 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END B2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.03 2.735 1.95 ;
        RECT 0.72 1.95 2.735 2.12 ;
        RECT 1.16 0.86 3.945 1.03 ;
        RECT 0.72 2.12 1.05 2.735 ;
        RECT 1.16 0.35 1.49 0.86 ;
        RECT 3.615 0.35 3.945 0.86 ;
    END
    ANTENNADIFFAREA 0.9326 ;
    ANTENNAPARTIALMETALSIDEAREA 1.361 LAYER li1 ;
  END Y

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.115 0.44 4.675 1.79 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.11 LAYER li1 ;
  END A1

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.26 3.82 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.103 LAYER li1 ;
  END B1

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.45 1.795 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END C1

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.895 1.45 1.295 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER li1 ;
  END D1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005 1.45 2.335 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END C2

  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.12 0.55 1.79 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.083 LAYER li1 ;
  END D2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.28 0.085 ;
      RECT 4.89 0.085 5.14 1.03 ;
      RECT 0.2 0.085 0.53 0.95 ;
      RECT 2.135 0.085 3.12 0.68 ;
      RECT 0 3.245 5.28 3.415 ;
      RECT 4.3 2.3 4.63 3.245 ;
      RECT 2.78 2.905 4.13 3.075 ;
      RECT 2.78 2.65 3.13 2.905 ;
      RECT 3.8 2.13 4.13 2.905 ;
      RECT 3.8 1.96 5.165 2.13 ;
      RECT 4.835 2.13 5.165 2.98 ;
      RECT 1.72 2.46 2.05 2.735 ;
      RECT 1.72 2.29 3.63 2.46 ;
      RECT 3.3 2.46 3.63 2.735 ;
      RECT 3.3 1.95 3.63 2.29 ;
      RECT 0.175 2.905 2.55 3.075 ;
      RECT 2.22 2.63 2.55 2.905 ;
      RECT 1.22 2.29 1.55 2.905 ;
      RECT 0.175 1.96 0.505 2.905 ;
    LAYER mcon ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_udb_a2222oi_1

MACRO scs8ls_udb_a2222oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.135 1.45 5.635 1.78 ;
        RECT 5.465 1.78 5.635 1.95 ;
        RECT 5.465 1.95 6.635 2.12 ;
        RECT 6.465 1.78 6.635 1.95 ;
        RECT 6.465 1.45 6.875 1.78 ;
    END
    ANTENNAGATEAREA 0.492 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.514 LAYER li1 ;
  END B1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.775 1.45 3.235 1.78 ;
        RECT 2.775 1.78 2.945 1.95 ;
        RECT 2.775 1.95 4.225 2.12 ;
        RECT 4.055 1.78 4.225 1.95 ;
        RECT 4.055 1.45 4.885 1.78 ;
    END
    ANTENNAGATEAREA 0.492 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.646 LAYER li1 ;
  END C2

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285 1.47 8.995 1.8 ;
        RECT 8.285 1.8 8.455 1.95 ;
        RECT 7.305 1.95 8.455 2.12 ;
        RECT 7.305 1.78 7.475 1.95 ;
        RECT 7.085 1.45 7.475 1.78 ;
    END
    ANTENNAGATEAREA 0.492 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.476 LAYER li1 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.705 1.45 8.035 1.78 ;
    END
    ANTENNAGATEAREA 0.492 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END A2

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.805 1.45 6.135 1.78 ;
    END
    ANTENNAGATEAREA 0.492 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405 1.45 3.735 1.78 ;
    END
    ANTENNAGATEAREA 0.492 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END C1

  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.42 1.45 2.275 1.78 ;
    END
    ANTENNAGATEAREA 0.492 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.101 LAYER li1 ;
  END D1

  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.255 0.935 0.67 ;
    END
    ANTENNAGATEAREA 0.492 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.081 LAYER li1 ;
  END D2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 0.81 5.26 1.11 ;
        RECT 1.08 1.11 8.99 1.28 ;
        RECT 4.93 0.35 5.26 0.81 ;
        RECT 1.08 1.28 1.25 1.94 ;
        RECT 1.635 1.025 1.965 1.11 ;
        RECT 3.52 0.595 3.69 1.11 ;
        RECT 6.85 0.35 7.18 1.11 ;
        RECT 8.66 0.35 8.99 1.11 ;
        RECT 0.92 1.94 1.25 1.95 ;
        RECT 0.92 1.95 2.4 2.12 ;
        RECT 0.92 2.12 1.25 2.735 ;
        RECT 2.07 2.12 2.4 2.735 ;
    END
    ANTENNADIFFAREA 1.9287 ;
    ANTENNAPARTIALMETALSIDEAREA 2.732 LAYER li1 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 5.44 0.77 6.68 0.94 ;
      RECT 5.44 0.35 5.69 0.77 ;
      RECT 6.43 0.35 6.68 0.77 ;
      RECT 7.35 0.77 8.48 0.94 ;
      RECT 7.35 0.35 7.6 0.77 ;
      RECT 8.31 0.35 8.48 0.77 ;
      RECT 3.01 0.255 4.2 0.425 ;
      RECT 3.87 0.425 4.2 0.94 ;
      RECT 3.01 0.425 3.34 0.94 ;
      RECT 1.135 0.855 1.465 0.94 ;
      RECT 1.135 0.605 2.44 0.855 ;
      RECT 2.57 2.29 4.725 2.46 ;
      RECT 4.395 2.46 4.725 2.735 ;
      RECT 4.395 1.95 4.725 2.29 ;
      RECT 0.42 2.905 2.9 3.075 ;
      RECT 2.57 2.46 2.9 2.905 ;
      RECT 0.42 1.94 0.75 2.905 ;
      RECT 1.57 2.29 1.9 2.905 ;
      RECT 3.945 2.96 6.635 3.075 ;
      RECT 3.1 2.905 6.635 2.96 ;
      RECT 3.1 2.63 4.195 2.905 ;
      RECT 5.485 2.63 5.655 2.905 ;
      RECT 6.385 2.63 6.635 2.905 ;
      RECT 4.955 2.29 9.005 2.46 ;
      RECT 8.675 2.46 9.005 2.98 ;
      RECT 5.855 2.46 6.185 2.735 ;
      RECT 6.805 2.46 7.135 2.98 ;
      RECT 6.805 1.95 7.135 2.29 ;
      RECT 4.955 2.46 5.285 2.735 ;
      RECT 4.955 1.95 5.285 2.29 ;
      RECT 0 -0.085 9.12 0.085 ;
      RECT 0.115 0.84 0.91 1.17 ;
      RECT 0.115 0.085 0.285 0.84 ;
      RECT 2.62 0.085 2.79 0.94 ;
      RECT 4.37 0.085 4.7 0.64 ;
      RECT 5.875 0.085 6.245 0.6 ;
      RECT 7.785 0.085 8.125 0.6 ;
      RECT 0 3.245 9.12 3.415 ;
      RECT 7.305 2.63 7.635 3.245 ;
      RECT 8.225 2.63 8.475 3.245 ;
    LAYER mcon ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
  END
END scs8ls_udb_a2222oi_2

MACRO scs8ls_udb_br0_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.96 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN DB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.35 0.875 2.92 ;
    END
    ANTENNADIFFAREA 0.1961 ;
    ANTENNAPARTIALMETALSIDEAREA 0.094 LAYER li1 ;
  END DB

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.35 0.425 2.18 ;
    END
    ANTENNAGATEAREA 0.111 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.092 LAYER li1 ;
  END EN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.96 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.96 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 0.96 3.415 ;
      RECT 0 -0.085 0.96 0.085 ;
      RECT 0.095 0.085 0.425 1.15 ;
    LAYER mcon ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_udb_br0_1

MACRO scs8ls_udb_br0_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN DB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.35 0.845 2.92 ;
    END
    ANTENNADIFFAREA 0.2072 ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER li1 ;
  END DB

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.35 0.425 2.18 ;
    END
    ANTENNAGATEAREA 0.222 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.092 LAYER li1 ;
  END EN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 1.44 3.415 ;
      RECT 0 -0.085 1.44 0.085 ;
      RECT 1.015 0.085 1.345 1.15 ;
      RECT 0.095 0.085 0.425 1.15 ;
    LAYER mcon ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_udb_br0_2

MACRO scs8ls_udb_bushold0_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN RESET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.525 1.355 2.195 ;
    END
    ANTENNAGATEAREA 0.126 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END RESET

  PIN X
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225 0.84 2.315 1.015 ;
        RECT 2.025 1.015 2.315 2.365 ;
        RECT 1.225 0.35 1.525 0.84 ;
        RECT 0.485 2.365 2.315 2.535 ;
        RECT 2.025 2.535 2.315 3.05 ;
        RECT 0.485 1.525 0.815 2.365 ;
    END
    ANTENNADIFFAREA 0.2289 ;
    ANTENNAGATEAREA 0.126 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.826 LAYER li1 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 2.4 3.415 ;
      RECT 0.815 2.72 1.145 3.245 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 1.975 0.085 2.305 0.61 ;
      RECT 0.795 0.085 1.055 0.69 ;
      RECT 0.085 1.185 1.855 1.355 ;
      RECT 1.605 1.355 1.855 2.195 ;
      RECT 0.085 2.72 0.425 3.05 ;
      RECT 0.085 1.355 0.315 2.72 ;
      RECT 0.085 1.055 0.625 1.185 ;
      RECT 0.335 0.35 0.625 1.055 ;
    LAYER mcon ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_udb_bushold0_1

MACRO scs8ls_udb_dec2to4_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.51 1.35 1.875 1.78 ;
        RECT 1.705 1.78 1.875 2.905 ;
        RECT 1.705 2.905 3.525 3.075 ;
        RECT 3.355 2.095 3.525 2.905 ;
        RECT 3.355 1.925 4.2 2.095 ;
        RECT 3.87 1.765 4.2 1.925 ;
    END
    ANTENNAGATEAREA 0.684 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.043 LAYER li1 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.705 1.625 ;
        RECT 0.535 0.705 0.705 1.18 ;
        RECT 0.535 0.59 3.44 0.705 ;
        RECT 1.485 0.705 3.44 0.76 ;
        RECT 0.535 0.535 1.655 0.59 ;
        RECT 3.27 0.76 3.44 1.425 ;
        RECT 3.27 1.425 4.12 1.595 ;
        RECT 3.27 1.595 3.63 1.755 ;
        RECT 3.95 0.71 4.12 1.425 ;
        RECT 3.95 0.54 6.025 0.71 ;
        RECT 5.855 0.71 6.025 1.01 ;
        RECT 5.855 1.01 6.775 1.18 ;
        RECT 6.445 1.18 6.775 1.55 ;
    END
    ANTENNAGATEAREA 0.684 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.035 LAYER li1 ;
  END A1

  PIN S1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.595 1.82 7.115 2.98 ;
        RECT 6.945 0.84 7.115 1.82 ;
        RECT 6.195 0.67 7.115 0.84 ;
        RECT 6.195 0.35 6.525 0.67 ;
    END
    ANTENNADIFFAREA 0.5376 ;
    ANTENNAPARTIALMETALSIDEAREA 0.576 LAYER li1 ;
  END S1

  PIN S0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.875 0.875 1.315 1.78 ;
        RECT 0.875 1.78 1.045 1.795 ;
        RECT 0.335 1.795 1.045 1.965 ;
        RECT 0.335 1.965 0.665 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
    ANTENNAPARTIALMETALSIDEAREA 0.481 LAYER li1 ;
  END S0

  PIN S3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.785 1.13 5.155 2.735 ;
        RECT 4.785 0.88 5.505 1.13 ;
    END
    ANTENNADIFFAREA 0.545 ;
    ANTENNAPARTIALMETALSIDEAREA 0.311 LAYER li1 ;
  END S3

  PIN S2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.18 2.56 2.735 ;
        RECT 1.815 0.93 2.23 1.18 ;
    END
    ANTENNADIFFAREA 0.5376 ;
    ANTENNAPARTIALMETALSIDEAREA 0.238 LAYER li1 ;
  END S2

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.73 2.265 3.185 2.725 ;
      RECT 2.73 0.93 3.1 2.265 ;
      RECT 0 -0.085 7.2 0.085 ;
      RECT 6.705 0.085 7.085 0.5 ;
      RECT 3.61 0.085 4.985 0.37 ;
      RECT 5.685 0.085 6.015 0.37 ;
      RECT 0.115 0.085 0.365 1.01 ;
      RECT 1.305 0.085 1.635 0.365 ;
      RECT 3.61 0.37 3.78 1.255 ;
      RECT 2.325 0.085 3.38 0.42 ;
      RECT 0 3.245 7.2 3.415 ;
      RECT 5.725 1.85 6.055 3.245 ;
      RECT 3.695 2.265 4.025 3.245 ;
      RECT 1.205 2.135 1.535 3.245 ;
      RECT 5.385 1.35 6.175 1.68 ;
      RECT 4.195 2.905 5.555 3.075 ;
      RECT 5.385 1.68 5.555 2.905 ;
      RECT 4.195 2.265 4.54 2.905 ;
      RECT 4.37 1.31 4.54 2.265 ;
      RECT 4.29 0.88 4.54 1.31 ;
    LAYER mcon ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_udb_dec2to4_1

MACRO scs8ls_udb_dlclkrn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.305 0.35 6.635 1.82 ;
        RECT 6.225 1.82 6.635 2.075 ;
    END
    ANTENNADIFFAREA 0.5376 ;
    ANTENNAPARTIALMETALSIDEAREA 0.155 LAYER li1 ;
  END GCLK

  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.845 1.29 7.225 1.96 ;
    END
    ANTENNAGATEAREA 0.516 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.142 LAYER li1 ;
  END CLKN

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.18 5.325 1.55 ;
    END
    ANTENNAGATEAREA 0.261 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.086 LAYER li1 ;
  END RESETB

  PIN GATEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955 1.445 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.071 LAYER li1 ;
  END GATEN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.995 1.915 2.69 2.245 ;
      RECT 2.52 1.02 2.69 1.915 ;
      RECT 2.52 0.85 4.24 1.02 ;
      RECT 3.925 1.02 4.24 1.655 ;
      RECT 1.65 0.48 3.05 0.85 ;
      RECT 0.085 1.105 2.35 1.275 ;
      RECT 2.035 1.275 2.35 1.745 ;
      RECT 2.035 1.075 2.35 1.105 ;
      RECT 0.085 2.29 0.56 2.795 ;
      RECT 0.085 1.275 0.255 2.29 ;
      RECT 0.085 0.35 0.51 1.105 ;
      RECT 3.385 1.825 5.865 2.075 ;
      RECT 5.535 1.225 5.865 1.825 ;
      RECT 3.385 1.3 3.715 1.825 ;
      RECT 4.41 0.35 4.66 1.825 ;
      RECT 2.86 2.245 7.565 2.415 ;
      RECT 7.235 2.415 7.565 2.98 ;
      RECT 7.235 2.13 7.565 2.245 ;
      RECT 7.395 1.12 7.565 2.13 ;
      RECT 7.235 0.35 7.565 1.12 ;
      RECT 1.495 2.415 3.03 2.585 ;
      RECT 1.495 2.12 1.825 2.415 ;
      RECT 2.86 1.235 3.175 2.245 ;
      RECT 0.425 1.95 1.825 2.12 ;
      RECT 1.495 1.445 1.825 1.95 ;
      RECT 0.425 1.445 0.745 1.95 ;
      RECT 0 -0.085 7.68 0.085 ;
      RECT 6.815 0.085 7.065 1.12 ;
      RECT 0.74 0.085 1.07 0.935 ;
      RECT 3.54 0.085 4.1 0.68 ;
      RECT 5.15 0.085 6.135 0.68 ;
      RECT 0 3.245 7.68 3.415 ;
      RECT 3.59 2.585 3.92 3.245 ;
      RECT 5.345 2.585 5.675 3.245 ;
      RECT 6.785 2.585 7.035 3.245 ;
      RECT 0.765 2.29 1.095 3.245 ;
    LAYER mcon ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
  END
END scs8ls_udb_dlclkrn_1

MACRO scs8ls_udb_dlclkrn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.67 0.81 7.525 1.01 ;
        RECT 5.67 1.01 6.595 1.13 ;
        RECT 5.67 0.35 6 0.81 ;
        RECT 7.195 0.35 7.525 0.81 ;
        RECT 6.365 1.13 6.595 1.865 ;
        RECT 6.365 1.865 7.065 2.035 ;
    END
    ANTENNADIFFAREA 0.8355 ;
    ANTENNAPARTIALMETALSIDEAREA 0.758 LAYER li1 ;
  END GCLK

  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.845 1.18 8.025 1.55 ;
    END
    ANTENNAGATEAREA 0.795 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.174 LAYER li1 ;
  END CLKN

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.18 5.305 1.55 ;
    END
    ANTENNAGATEAREA 0.261 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.082 LAYER li1 ;
  END RESETB

  PIN GATEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935 1.445 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.075 LAYER li1 ;
  END GATEN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 5.215 2.715 5.545 2.945 ;
      RECT 5.215 2.545 7.515 2.715 ;
      RECT 6.285 2.715 6.615 2.945 ;
      RECT 7.185 2.715 7.515 2.945 ;
      RECT 5.215 2.4 5.545 2.545 ;
      RECT 1.825 2.405 2.665 2.735 ;
      RECT 2.495 1.02 2.665 2.405 ;
      RECT 2.495 0.85 4.22 1.02 ;
      RECT 3.89 1.02 4.22 1.335 ;
      RECT 1.63 0.48 2.835 0.85 ;
      RECT 0.085 1.105 2.325 1.275 ;
      RECT 2.025 1.275 2.325 1.775 ;
      RECT 0.085 2.29 0.575 2.795 ;
      RECT 0.085 1.275 0.255 2.29 ;
      RECT 0.255 0.35 0.6 1.105 ;
      RECT 3.35 1.72 5.685 1.89 ;
      RECT 5.515 1.645 5.685 1.72 ;
      RECT 5.515 1.315 6.185 1.645 ;
      RECT 4.07 1.89 4.4 2.03 ;
      RECT 3.35 1.31 3.68 1.72 ;
      RECT 4.39 0.35 4.64 1.72 ;
      RECT 2.835 2.205 7.405 2.23 ;
      RECT 5.715 2.23 7.405 2.375 ;
      RECT 7.235 1.93 7.405 2.205 ;
      RECT 7.235 1.76 8.525 1.93 ;
      RECT 8.195 1.93 8.525 2.98 ;
      RECT 8.195 0.35 8.525 1.76 ;
      RECT 2.835 2.2 5.885 2.205 ;
      RECT 4.57 2.06 5.885 2.2 ;
      RECT 1.485 2.905 3.14 3.075 ;
      RECT 2.835 2.37 3.14 2.905 ;
      RECT 1.485 2.12 1.655 2.905 ;
      RECT 2.835 2.23 4.74 2.37 ;
      RECT 0.425 1.95 1.655 2.12 ;
      RECT 1.485 1.775 1.655 1.95 ;
      RECT 1.485 1.445 1.815 1.775 ;
      RECT 2.835 1.26 3.14 2.2 ;
      RECT 0.425 1.445 0.725 1.95 ;
      RECT 0 -0.085 8.64 0.085 ;
      RECT 7.695 0.085 8.025 1.01 ;
      RECT 0.77 0.085 1.1 0.935 ;
      RECT 3.325 0.085 4.08 0.68 ;
      RECT 5.13 0.085 5.46 1.01 ;
      RECT 6.17 0.085 7.025 0.6 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 5.75 2.885 6.08 3.245 ;
      RECT 3.53 2.54 3.865 3.245 ;
      RECT 4.605 2.54 4.985 3.245 ;
      RECT 0.785 2.29 1.115 3.245 ;
      RECT 7.745 2.1 7.995 3.245 ;
    LAYER mcon ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
  END
END scs8ls_udb_dlclkrn_2

MACRO scs8ls_udb_dlclkrn_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.56 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.325 1.39 8.085 1.78 ;
        RECT 7.755 1.78 8.085 1.82 ;
        RECT 6.765 1.22 8.095 1.39 ;
        RECT 7.755 1.82 8.985 2.07 ;
        RECT 6.765 1.13 7.095 1.22 ;
        RECT 7.765 1.01 8.095 1.22 ;
        RECT 5.71 0.96 7.095 1.13 ;
        RECT 7.765 0.84 9.095 1.01 ;
        RECT 5.71 0.35 6.04 0.96 ;
        RECT 6.765 0.35 7.095 0.96 ;
        RECT 7.765 0.35 8.095 0.84 ;
        RECT 8.765 0.35 9.095 0.84 ;
    END
    ANTENNADIFFAREA 1.5378 ;
    ANTENNAPARTIALMETALSIDEAREA 1.459 LAYER li1 ;
  END GCLK

  PIN GATEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.45 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1 ;
  END GATEN

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.18 5.345 1.54 ;
    END
    ANTENNAGATEAREA 0.279 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER li1 ;
  END RESETB

  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 8.285 1.18 9.475 1.55 ;
    END
    ANTENNAGATEAREA 1.353 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.108 LAYER li1 ;
  END CLKN

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.56 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.56 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.825 2.07 2.715 2.4 ;
      RECT 2.545 1.09 2.715 2.07 ;
      RECT 2.545 0.92 4.295 1.09 ;
      RECT 3.965 1.09 4.295 1.54 ;
      RECT 1.66 0.48 2.83 0.92 ;
      RECT 3.425 1.71 5.725 1.88 ;
      RECT 5.555 1.63 5.725 1.71 ;
      RECT 5.555 1.3 6.595 1.63 ;
      RECT 4.145 1.88 4.555 2.11 ;
      RECT 3.425 1.31 3.755 1.71 ;
      RECT 4.48 0.75 4.65 1.71 ;
      RECT 4.32 0.35 4.65 0.75 ;
      RECT 0.085 1.1 2.375 1.27 ;
      RECT 2.045 1.27 2.375 1.79 ;
      RECT 0.085 1.94 0.455 2.82 ;
      RECT 0.085 1.27 0.255 1.94 ;
      RECT 0.085 0.35 0.59 1.1 ;
      RECT 6.735 2.24 9.495 2.41 ;
      RECT 9.325 1.93 9.495 2.24 ;
      RECT 9.325 1.76 10.255 1.93 ;
      RECT 10.085 1.93 10.255 2.1 ;
      RECT 9.765 0.35 10.255 1.76 ;
      RECT 10.085 2.1 10.445 2.98 ;
      RECT 2.885 2.28 5.065 2.45 ;
      RECT 4.895 2.22 5.065 2.28 ;
      RECT 4.895 2.05 6.065 2.22 ;
      RECT 5.895 1.97 6.065 2.05 ;
      RECT 5.895 1.8 6.905 1.97 ;
      RECT 6.735 1.97 6.905 2.24 ;
      RECT 1.485 2.57 3.215 2.74 ;
      RECT 2.885 2.45 3.215 2.57 ;
      RECT 1.485 2.12 1.655 2.57 ;
      RECT 0.625 1.95 1.655 2.12 ;
      RECT 2.885 1.26 3.215 2.28 ;
      RECT 1.485 1.8 1.655 1.95 ;
      RECT 1.485 1.47 1.835 1.8 ;
      RECT 0.625 1.77 0.795 1.95 ;
      RECT 0.425 1.44 0.795 1.77 ;
      RECT 6.235 2.75 6.565 2.98 ;
      RECT 6.235 2.58 9.435 2.75 ;
      RECT 7.305 2.75 7.635 2.98 ;
      RECT 8.205 2.75 8.535 2.98 ;
      RECT 9.105 2.75 9.435 2.98 ;
      RECT 6.235 2.56 6.565 2.58 ;
      RECT 5.235 2.39 6.565 2.56 ;
      RECT 5.235 2.56 5.565 2.98 ;
      RECT 6.235 2.14 6.565 2.39 ;
      RECT 0 -0.085 10.56 0.085 ;
      RECT 9.265 0.085 9.595 1.01 ;
      RECT 0.76 0.085 1.09 0.93 ;
      RECT 3.4 0.085 4.09 0.68 ;
      RECT 5.14 0.085 5.47 1.01 ;
      RECT 6.21 0.085 6.54 0.79 ;
      RECT 7.265 0.085 7.595 1.05 ;
      RECT 8.265 0.085 8.595 0.67 ;
      RECT 0 3.245 10.56 3.415 ;
      RECT 6.77 2.92 7.1 3.245 ;
      RECT 5.735 2.73 6.065 3.245 ;
      RECT 3.63 2.62 4.025 3.245 ;
      RECT 4.675 2.62 5.005 3.245 ;
      RECT 0.785 2.29 1.115 3.245 ;
      RECT 9.665 2.1 9.915 3.245 ;
    LAYER mcon ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_udb_dlclkrn_4

MACRO scs8ls_udb_dlclkrp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.195 1.82 8.555 2.98 ;
        RECT 8.385 1.13 8.555 1.82 ;
        RECT 8.275 0.35 8.555 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
    ANTENNAPARTIALMETALSIDEAREA 0.416 LAYER li1 ;
  END GCLK

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.32 1.18 6.65 1.55 ;
    END
    ANTENNAGATEAREA 0.498 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.072 LAYER li1 ;
  END CLK

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.26 1.35 4.675 2.02 ;
    END
    ANTENNAGATEAREA 0.222 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.149 LAYER li1 ;
  END RESETB

  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.99 1.545 1.77 1.8 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.071 LAYER li1 ;
  END GATE

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.09 1.97 2.79 2.14 ;
      RECT 2.52 1.47 2.79 1.97 ;
      RECT 0.09 2.14 0.52 2.82 ;
      RECT 0.09 1.94 0.57 1.97 ;
      RECT 0.09 1.035 0.26 1.94 ;
      RECT 0.09 0.35 0.545 1.035 ;
      RECT 7.855 1.3 8.215 1.63 ;
      RECT 7.16 1.97 7.49 2.86 ;
      RECT 7.16 1.8 8.025 1.97 ;
      RECT 7.855 1.63 8.025 1.8 ;
      RECT 7.855 1.13 8.025 1.3 ;
      RECT 7.205 0.96 8.025 1.13 ;
      RECT 7.205 0.35 7.535 0.96 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 4.04 2.53 4.21 3.245 ;
      RECT 4.97 2.53 5.3 3.245 ;
      RECT 0.69 2.31 1.62 3.245 ;
      RECT 7.695 2.14 8.025 3.245 ;
      RECT 6.74 2.06 6.99 3.245 ;
      RECT 0 -0.085 8.64 0.085 ;
      RECT 0.715 0.085 1.045 1.03 ;
      RECT 3.7 0.085 4.75 0.5 ;
      RECT 6.385 0.085 6.715 1.01 ;
      RECT 7.765 0.085 8.095 0.79 ;
      RECT 5.47 2.87 6.57 3.04 ;
      RECT 6.4 1.89 6.57 2.87 ;
      RECT 6.4 1.72 6.99 1.89 ;
      RECT 6.82 1.63 6.99 1.72 ;
      RECT 6.82 1.3 7.68 1.63 ;
      RECT 5.47 1.82 5.75 2.87 ;
      RECT 5.47 1.18 5.64 1.82 ;
      RECT 3.7 1.01 5.64 1.18 ;
      RECT 5.26 0.595 5.64 1.01 ;
      RECT 3.7 1.18 4.03 1.805 ;
      RECT 3.36 0.67 5.09 0.84 ;
      RECT 4.92 0.425 5.09 0.67 ;
      RECT 4.92 0.255 6.15 0.425 ;
      RECT 5.82 0.425 6.15 1.13 ;
      RECT 5.98 1.13 6.15 1.82 ;
      RECT 5.98 1.82 6.23 2.7 ;
      RECT 3.3 2.045 3.53 2.375 ;
      RECT 3.36 0.84 3.53 2.045 ;
      RECT 3.36 0.45 3.53 0.67 ;
      RECT 1.53 0.28 3.53 0.45 ;
      RECT 1.53 0.45 1.74 1.205 ;
      RECT 0.43 1.205 2.31 1.375 ;
      RECT 1.98 1.375 2.31 1.8 ;
      RECT 0.43 1.375 0.75 1.605 ;
      RECT 3.7 2.19 5.015 2.36 ;
      RECT 4.41 2.36 4.74 2.975 ;
      RECT 4.845 1.68 5.015 2.19 ;
      RECT 4.845 1.35 5.3 1.68 ;
      RECT 2.675 2.545 3.87 2.875 ;
      RECT 3.7 2.36 3.87 2.545 ;
      RECT 2.96 0.95 3.13 2.545 ;
      RECT 2.105 0.62 3.13 0.95 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_udb_dlclkrp_1

MACRO scs8ls_udb_dlclkrp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.195 1.82 8.535 2.98 ;
        RECT 8.365 1.13 8.535 1.82 ;
        RECT 8.275 0.35 8.535 1.13 ;
    END
    ANTENNADIFFAREA 0.5432 ;
    ANTENNAPARTIALMETALSIDEAREA 0.408 LAYER li1 ;
  END GCLK

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.32 1.18 6.65 1.55 ;
    END
    ANTENNAGATEAREA 0.498 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.072 LAYER li1 ;
  END CLK

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.26 1.35 4.675 2.02 ;
    END
    ANTENNAGATEAREA 0.222 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.149 LAYER li1 ;
  END RESETB

  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.99 1.545 1.77 1.8 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.071 LAYER li1 ;
  END GATE

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.7 2.19 5.015 2.36 ;
      RECT 4.41 2.36 4.74 2.975 ;
      RECT 4.845 1.68 5.015 2.19 ;
      RECT 4.845 1.35 5.3 1.68 ;
      RECT 2.665 2.545 3.87 2.875 ;
      RECT 3.7 2.36 3.87 2.545 ;
      RECT 2.96 0.95 3.13 2.545 ;
      RECT 2.105 0.62 3.13 0.95 ;
      RECT 0.09 1.97 2.79 2.14 ;
      RECT 2.52 1.47 2.79 1.97 ;
      RECT 0.09 2.14 0.52 2.82 ;
      RECT 0.09 1.94 0.57 1.97 ;
      RECT 0.09 1.035 0.26 1.94 ;
      RECT 0.09 0.35 0.545 1.035 ;
      RECT 0 3.245 9.12 3.415 ;
      RECT 8.71 1.82 8.975 3.245 ;
      RECT 4.97 2.53 5.3 3.245 ;
      RECT 7.695 2.14 8.025 3.245 ;
      RECT 6.74 2.06 6.99 3.245 ;
      RECT 4.04 2.53 4.21 3.245 ;
      RECT 0.69 2.31 1.62 3.245 ;
      RECT 5.47 2.87 6.57 3.04 ;
      RECT 6.4 1.89 6.57 2.87 ;
      RECT 6.4 1.72 6.99 1.89 ;
      RECT 6.82 1.63 6.99 1.72 ;
      RECT 6.82 1.3 7.68 1.63 ;
      RECT 5.47 1.82 5.75 2.87 ;
      RECT 5.47 1.18 5.64 1.82 ;
      RECT 3.7 1.01 5.64 1.18 ;
      RECT 5.26 0.595 5.64 1.01 ;
      RECT 3.7 1.18 4.03 1.805 ;
      RECT 7.16 1.97 7.49 2.86 ;
      RECT 7.16 1.8 8.025 1.97 ;
      RECT 7.855 1.63 8.025 1.8 ;
      RECT 7.855 1.3 8.195 1.63 ;
      RECT 7.855 1.13 8.025 1.3 ;
      RECT 7.205 0.96 8.025 1.13 ;
      RECT 7.205 0.35 7.535 0.96 ;
      RECT 0 -0.085 9.12 0.085 ;
      RECT 8.705 0.085 8.955 1.13 ;
      RECT 0.715 0.085 1.045 1.03 ;
      RECT 3.7 0.085 4.75 0.5 ;
      RECT 6.385 0.085 6.715 1.01 ;
      RECT 7.765 0.085 8.095 0.79 ;
      RECT 3.36 0.67 5.09 0.84 ;
      RECT 4.92 0.425 5.09 0.67 ;
      RECT 4.92 0.255 6.15 0.425 ;
      RECT 5.82 0.425 6.15 1.13 ;
      RECT 5.98 1.13 6.15 1.82 ;
      RECT 5.98 1.82 6.23 2.7 ;
      RECT 3.3 2.045 3.53 2.375 ;
      RECT 3.36 0.84 3.53 2.045 ;
      RECT 3.36 0.45 3.53 0.67 ;
      RECT 1.53 0.28 3.53 0.45 ;
      RECT 1.53 0.45 1.74 1.205 ;
      RECT 0.43 1.205 2.31 1.375 ;
      RECT 1.98 1.375 2.31 1.8 ;
      RECT 0.43 1.375 0.75 1.605 ;
    LAYER mcon ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_udb_dlclkrp_2

MACRO scs8ls_udb_dlclkrp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 10.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.195 1.975 8.535 2.98 ;
        RECT 8.195 1.805 9.465 1.975 ;
        RECT 9.13 1.975 9.465 2.98 ;
        RECT 9.13 1.325 9.465 1.805 ;
        RECT 9.13 1.13 9.36 1.325 ;
        RECT 8.275 0.96 9.36 1.13 ;
        RECT 8.275 0.35 8.45 0.96 ;
        RECT 9.13 0.35 9.36 0.96 ;
    END
    ANTENNADIFFAREA 1.0864 ;
    ANTENNAPARTIALMETALSIDEAREA 0.798 LAYER li1 ;
  END GCLK

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.32 1.18 6.65 1.55 ;
    END
    ANTENNAGATEAREA 0.498 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.072 LAYER li1 ;
  END CLK

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.26 1.35 4.675 2.02 ;
    END
    ANTENNAGATEAREA 0.222 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.149 LAYER li1 ;
  END RESETB

  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.99 1.545 1.77 1.8 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.071 LAYER li1 ;
  END GATE

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 10.08 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 10.08 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.36 0.67 5.09 0.84 ;
      RECT 4.92 0.425 5.09 0.67 ;
      RECT 4.92 0.255 6.15 0.425 ;
      RECT 5.82 0.425 6.15 1.13 ;
      RECT 5.98 1.13 6.15 1.82 ;
      RECT 5.98 1.82 6.23 2.7 ;
      RECT 3.3 2.045 3.53 2.375 ;
      RECT 3.36 0.84 3.53 2.045 ;
      RECT 3.36 0.45 3.53 0.67 ;
      RECT 1.53 0.28 3.53 0.45 ;
      RECT 1.53 0.45 1.74 1.205 ;
      RECT 0.43 1.205 2.31 1.375 ;
      RECT 1.98 1.375 2.31 1.8 ;
      RECT 0.43 1.375 0.75 1.605 ;
      RECT 7.855 1.3 8.9 1.63 ;
      RECT 7.16 1.97 7.49 2.86 ;
      RECT 7.16 1.8 8.025 1.97 ;
      RECT 7.855 1.63 8.025 1.8 ;
      RECT 7.855 1.13 8.025 1.3 ;
      RECT 7.205 0.96 8.025 1.13 ;
      RECT 7.205 0.35 7.535 0.96 ;
      RECT 0 -0.085 10.08 0.085 ;
      RECT 9.53 0.085 9.815 1.13 ;
      RECT 0.715 0.085 1.045 1.03 ;
      RECT 3.7 0.085 4.75 0.5 ;
      RECT 6.385 0.085 6.715 1.01 ;
      RECT 7.765 0.085 8.095 0.79 ;
      RECT 8.625 0.085 8.955 0.79 ;
      RECT 3.7 2.19 5.015 2.36 ;
      RECT 4.41 2.36 4.74 2.975 ;
      RECT 4.845 1.68 5.015 2.19 ;
      RECT 4.845 1.35 5.3 1.68 ;
      RECT 2.665 2.545 3.87 2.875 ;
      RECT 3.7 2.36 3.87 2.545 ;
      RECT 2.96 0.95 3.13 2.545 ;
      RECT 2.105 0.62 3.13 0.95 ;
      RECT 0.09 1.97 2.79 2.14 ;
      RECT 2.52 1.47 2.79 1.97 ;
      RECT 0.09 2.14 0.52 2.82 ;
      RECT 0.09 1.94 0.57 1.97 ;
      RECT 0.09 1.035 0.26 1.94 ;
      RECT 0.09 0.35 0.545 1.035 ;
      RECT 0 3.245 10.08 3.415 ;
      RECT 9.635 1.82 9.885 3.245 ;
      RECT 4.97 2.53 5.3 3.245 ;
      RECT 7.695 2.14 8.025 3.245 ;
      RECT 6.74 2.06 6.99 3.245 ;
      RECT 8.705 2.15 8.96 3.245 ;
      RECT 4.04 2.53 4.21 3.245 ;
      RECT 0.69 2.31 1.62 3.245 ;
      RECT 5.47 2.87 6.57 3.04 ;
      RECT 6.4 1.89 6.57 2.87 ;
      RECT 6.4 1.72 6.99 1.89 ;
      RECT 6.82 1.63 6.99 1.72 ;
      RECT 6.82 1.3 7.68 1.63 ;
      RECT 5.47 1.82 5.75 2.87 ;
      RECT 5.47 1.18 5.64 1.82 ;
      RECT 3.7 1.01 5.64 1.18 ;
      RECT 5.26 0.595 5.64 1.01 ;
      RECT 3.7 1.18 4.03 1.805 ;
    LAYER mcon ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_udb_dlclkrp_4

MACRO scs8ls_udb_emux2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.515 1.45 7.075 1.78 ;
    END
    ANTENNAGATEAREA 0.261 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.11 LAYER li1 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.245 1.3 7.575 1.78 ;
    END
    ANTENNAGATEAREA 0.261 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.094 LAYER li1 ;
  END A1

  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.95 1.45 5.35 1.78 ;
    END
    ANTENNAGATEAREA 0.4695 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER li1 ;
  END S

  PIN TEB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.35 3.6 1.68 ;
        RECT 1.565 1.68 3.235 1.72 ;
        RECT 0.425 1.72 3.235 1.89 ;
        RECT 0.425 1.56 0.755 1.72 ;
    END
    ANTENNAGATEAREA 0.5445 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.503 LAYER li1 ;
  END TEB

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 0.4 3.56 0.67 ;
        RECT 3.39 0.67 3.56 1.01 ;
        RECT 3.39 1.01 3.94 1.18 ;
        RECT 3.77 1.18 3.94 2.06 ;
        RECT 1.655 2.06 3.94 2.23 ;
        RECT 1.655 2.23 1.985 2.31 ;
    END
    ANTENNADIFFAREA 0.5432 ;
    ANTENNAPARTIALMETALSIDEAREA 0.98 LAYER li1 ;
  END Z

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 4.745 2.51 5.075 2.98 ;
      RECT 4.745 2.34 6.635 2.51 ;
      RECT 6.305 2.51 6.635 2.735 ;
      RECT 4.745 2.29 5.075 2.34 ;
      RECT 5.745 2.905 7.565 3.075 ;
      RECT 5.745 2.68 6.075 2.905 ;
      RECT 7.235 2.34 7.565 2.905 ;
      RECT 6.175 2 7.115 2.17 ;
      RECT 4.61 1.11 6.99 1.28 ;
      RECT 6.66 0.595 6.99 1.11 ;
      RECT 6.175 1.28 6.345 2 ;
      RECT 4.61 1.28 4.78 1.32 ;
      RECT 4.45 1.32 4.78 1.65 ;
      RECT 0.085 1.22 1.295 1.39 ;
      RECT 0.965 1.39 1.295 1.55 ;
      RECT 0.085 0.54 0.48 1.22 ;
      RECT 0.085 2.1 0.365 2.98 ;
      RECT 0.085 1.39 0.255 2.1 ;
      RECT 2.11 1.05 3.22 1.18 ;
      RECT 1.09 0.88 3.22 1.05 ;
      RECT 2.11 0.84 3.22 0.88 ;
      RECT 1.09 0.35 1.34 0.88 ;
      RECT 1.155 2.57 2.435 2.65 ;
      RECT 2.105 2.65 2.435 2.98 ;
      RECT 1.155 2.48 3.53 2.57 ;
      RECT 3.2 2.57 3.53 2.98 ;
      RECT 2.265 2.4 3.53 2.48 ;
      RECT 1.155 2.65 1.485 2.98 ;
      RECT 1.155 2.06 1.485 2.48 ;
      RECT 4.11 1.95 5.765 2.12 ;
      RECT 5.595 1.8 5.765 1.95 ;
      RECT 5.595 1.47 5.925 1.8 ;
      RECT 4.11 2.12 4.515 2.7 ;
      RECT 4.11 1.82 4.515 1.95 ;
      RECT 4.11 1.15 4.28 1.82 ;
      RECT 4.11 0.605 4.44 1.15 ;
      RECT 4.78 0.77 6.49 0.94 ;
      RECT 6.32 0.425 6.49 0.77 ;
      RECT 4.78 0.35 5.11 0.77 ;
      RECT 6.32 0.255 7.54 0.425 ;
      RECT 7.21 0.425 7.54 1.13 ;
      RECT 0 -0.085 7.68 0.085 ;
      RECT 3.73 0.085 3.93 0.84 ;
      RECT 5.28 0.085 6.15 0.6 ;
      RECT 0.66 0.085 0.91 1.05 ;
      RECT 1.52 0.085 1.85 0.71 ;
      RECT 0 3.245 7.68 3.415 ;
      RECT 2.665 2.74 2.995 3.245 ;
      RECT 5.245 2.68 5.575 3.245 ;
      RECT 3.73 2.4 3.9 3.245 ;
      RECT 0.565 2.1 0.895 3.245 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
  END
END scs8ls_udb_emux2_2

MACRO scs8ls_udb_fasumb_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.8 2.755 2.15 ;
        RECT 1.735 1.47 2.755 1.8 ;
    END
    ANTENNAGATEAREA 0.804 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.842 LAYER met1 ;
  END CIN

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.765 1.35 7.095 1.78 ;
    END
    ANTENNAGATEAREA 1.05 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 4.858 LAYER met1 ;
  END A

  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.43 0.39 8.035 1.17 ;
        RECT 7.805 1.17 8.035 1.84 ;
        RECT 7.605 1.84 8.035 2.98 ;
    END
    ANTENNADIFFAREA 0.5413 ;
    ANTENNAPARTIALMETALSIDEAREA 0.203 LAYER li1 ;
  END COUT

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525 0.92 6.255 1.09 ;
        RECT 2.525 0.81 3.235 0.92 ;
        RECT 4.275 1.09 4.605 1.59 ;
        RECT 5.925 1.09 6.255 1.59 ;
        RECT 2.525 0.425 2.695 0.81 ;
        RECT 1.13 0.255 2.695 0.425 ;
        RECT 1.13 0.425 1.46 0.57 ;
    END
    ANTENNAGATEAREA 1.05 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.285 LAYER li1 ;
  END B

  PIN SUMB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.94 0.42 6.595 0.75 ;
        RECT 6.425 0.75 6.595 2.32 ;
        RECT 5.315 2.32 6.595 2.49 ;
        RECT 5.315 2.49 5.565 2.735 ;
    END
    ANTENNADIFFAREA 1.0376 ;
    ANTENNAPARTIALMETALSIDEAREA 0.948 LAYER li1 ;
  END SUMB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.16 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 0.575 1.735 0.865 1.78 ;
      RECT 0.575 1.595 7.105 1.735 ;
      RECT 2.975 1.735 3.265 1.78 ;
      RECT 6.815 1.735 7.105 1.78 ;
      RECT 0.575 1.55 0.865 1.595 ;
      RECT 2.975 1.55 3.265 1.595 ;
      RECT 6.815 1.55 7.105 1.595 ;
      RECT 2.015 2.105 2.305 2.15 ;
      RECT 2.015 1.965 5.665 2.105 ;
      RECT 3.455 2.105 3.745 2.15 ;
      RECT 5.375 2.105 5.665 2.15 ;
      RECT 2.015 1.92 2.305 1.965 ;
      RECT 3.455 1.92 3.745 1.965 ;
      RECT 5.375 1.92 5.665 1.965 ;
    LAYER li1 ;
      RECT 7.265 1.34 7.635 1.67 ;
      RECT 4.975 2.905 6.935 3.075 ;
      RECT 6.765 2.12 6.935 2.905 ;
      RECT 6.765 1.95 7.435 2.12 ;
      RECT 7.265 1.67 7.435 1.95 ;
      RECT 1.975 2.8 2.305 2.98 ;
      RECT 1.975 2.49 2.305 2.63 ;
      RECT 1.565 2.32 2.305 2.49 ;
      RECT 1.395 1.08 2.25 1.25 ;
      RECT 1.92 0.66 2.25 1.08 ;
      RECT 1.395 1.25 1.565 1.97 ;
      RECT 1.565 2.14 1.735 2.32 ;
      RECT 1.395 1.97 1.735 2.14 ;
      RECT 1.975 2.63 5.145 2.8 ;
      RECT 4.975 2.8 5.145 2.905 ;
      RECT 4.975 1.65 5.145 2.63 ;
      RECT 4.815 1.32 5.145 1.65 ;
      RECT 0 3.245 8.16 3.415 ;
      RECT 7.105 2.29 7.435 3.245 ;
      RECT 2.93 2.97 3.26 3.245 ;
      RECT 4 2.97 4.35 3.245 ;
      RECT 0.615 2.65 1.055 3.245 ;
      RECT 0 -0.085 8.16 0.085 ;
      RECT 6.765 0.085 7.095 1.17 ;
      RECT 0.555 0.085 0.885 0.96 ;
      RECT 2.9 0.085 3.235 0.64 ;
      RECT 3.915 0.085 4.26 0.41 ;
      RECT 0.22 1.47 0.89 1.8 ;
      RECT 0.125 1.13 1.225 1.3 ;
      RECT 1.055 0.91 1.225 1.13 ;
      RECT 0.125 0.66 0.375 1.13 ;
      RECT 1.055 0.74 1.74 0.91 ;
      RECT 1.225 2.66 1.805 2.91 ;
      RECT 1.225 2.48 1.395 2.66 ;
      RECT 0.115 2.31 1.395 2.48 ;
      RECT 0.115 2.48 0.445 2.98 ;
      RECT 0.115 1.97 0.445 2.31 ;
      RECT 2.985 1.59 3.235 1.78 ;
      RECT 2.985 1.26 3.315 1.59 ;
      RECT 3.485 1.35 4.035 2.12 ;
      RECT 3.405 0.58 4.77 0.75 ;
      RECT 3.405 0.39 3.735 0.58 ;
      RECT 4.44 0.39 4.77 0.58 ;
      RECT 3.465 2.29 4.805 2.46 ;
      RECT 4.555 1.82 4.805 2.29 ;
      RECT 5.385 1.35 5.715 2.15 ;
    LAYER mcon ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.875 1.58 7.045 1.75 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 1.95 5.605 2.12 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 1.95 3.685 2.12 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 1.58 3.205 1.75 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 1.95 2.245 2.12 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 1.58 0.805 1.75 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_udb_fasumb_1

MACRO scs8ls_udb_mux3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.45 6.81 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.087 LAYER li1 ;
  END A0

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.05 1.45 7.555 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.099 LAYER li1 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.435 1.465 1.78 ;
    END
    ANTENNAGATEAREA 0.246 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.077 LAYER li1 ;
  END A2

  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.445 3.335 1.78 ;
    END
    ANTENNAGATEAREA 0.492 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.065 LAYER li1 ;
  END S1

  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925 1.45 5.255 1.78 ;
    END
    ANTENNAGATEAREA 0.492 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END S0

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.82 0.575 2.98 ;
        RECT 0.085 1.13 0.255 1.82 ;
        RECT 0.085 0.35 0.41 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
    ANTENNAPARTIALMETALSIDEAREA 0.451 LAYER li1 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 4.765 2.905 6.655 3.075 ;
      RECT 4.765 2.685 5.095 2.905 ;
      RECT 6.325 2.63 6.655 2.905 ;
      RECT 5.765 2.46 6.095 2.735 ;
      RECT 5.765 2.29 7.565 2.46 ;
      RECT 7.235 2.46 7.565 2.98 ;
      RECT 7.235 1.95 7.565 2.29 ;
      RECT 1.09 0.765 1.42 0.925 ;
      RECT 1.09 0.595 2.975 0.765 ;
      RECT 2.67 0.765 2.975 0.925 ;
      RECT 1.09 0.45 1.42 0.595 ;
      RECT 4.585 1.11 5.825 1.28 ;
      RECT 5.495 1.28 5.825 1.775 ;
      RECT 4.585 0.595 4.925 1.11 ;
      RECT 4.205 1.925 4.755 2.175 ;
      RECT 4.585 1.28 4.755 1.925 ;
      RECT 1.825 2.905 3.585 3.075 ;
      RECT 3.255 2.12 3.585 2.905 ;
      RECT 3.255 1.95 3.675 2.12 ;
      RECT 3.505 1.275 3.675 1.95 ;
      RECT 3.485 0.595 3.735 1.275 ;
      RECT 1.825 1.77 1.995 2.905 ;
      RECT 1.825 1.44 2.155 1.77 ;
      RECT 2.165 1.94 2.495 2.735 ;
      RECT 2.325 1.265 2.495 1.94 ;
      RECT 0.585 1.095 2.495 1.265 ;
      RECT 2.24 0.935 2.495 1.095 ;
      RECT 0.585 1.265 0.755 1.3 ;
      RECT 0.425 1.3 0.755 1.63 ;
      RECT 6.335 1.11 7.505 1.28 ;
      RECT 6.335 0.425 6.505 1.11 ;
      RECT 7.175 0.35 7.505 1.11 ;
      RECT 5.285 0.255 6.505 0.425 ;
      RECT 5.285 0.425 5.615 0.94 ;
      RECT 5.265 2.515 5.595 2.735 ;
      RECT 3.865 2.345 5.595 2.515 ;
      RECT 5.265 2.12 5.595 2.345 ;
      RECT 5.265 1.95 6.165 2.12 ;
      RECT 5.995 0.94 6.165 1.95 ;
      RECT 5.785 0.595 6.165 0.94 ;
      RECT 3.865 1.615 4.035 2.345 ;
      RECT 3.865 1.445 4.075 1.615 ;
      RECT 3.905 0.425 4.075 1.445 ;
      RECT 1.65 0.255 4.075 0.425 ;
      RECT 3.145 0.425 3.315 1.105 ;
      RECT 2.665 1.105 3.315 1.275 ;
      RECT 2.665 1.95 3.025 2.735 ;
      RECT 2.665 1.275 2.835 1.95 ;
      RECT 0.59 0.085 0.92 0.925 ;
      RECT 0 -0.085 7.68 0.085 ;
      RECT 4.245 0.085 4.415 1.275 ;
      RECT 6.675 0.085 7.005 0.94 ;
      RECT 0 3.245 7.68 3.415 ;
      RECT 3.755 2.685 4.085 3.245 ;
      RECT 6.855 2.65 7.035 3.245 ;
      RECT 0.745 1.95 1.075 3.245 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
  END
END scs8ls_udb_mux3_1

MACRO scs8ls_udb_srlb_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625 1.95 3.255 2.12 ;
        RECT 2.765 2.12 3.255 2.98 ;
        RECT 2.765 1.82 3.255 1.95 ;
        RECT 0.625 1.68 0.795 1.95 ;
        RECT 3.085 1.13 3.255 1.82 ;
        RECT 0.425 1.35 0.795 1.68 ;
        RECT 2.915 0.84 3.255 1.13 ;
        RECT 1.74 0.67 3.255 0.84 ;
        RECT 1.74 0.35 2.07 0.67 ;
        RECT 2.915 0.35 3.255 0.67 ;
    END
    ANTENNADIFFAREA 0.7707 ;
    ANTENNAGATEAREA 0.279 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.341 LAYER li1 ;
  END Q

  PIN R1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.35 1.835 1.78 ;
    END
    ANTENNAGATEAREA 0.279 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER li1 ;
  END R1

  PIN R2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.35 2.375 1.78 ;
    END
    ANTENNAGATEAREA 0.279 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER li1 ;
  END R2

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.85 0.455 2.98 ;
        RECT 0.085 1.18 0.255 1.85 ;
        RECT 0.085 1.01 2.745 1.18 ;
        RECT 2.575 1.18 2.745 1.3 ;
        RECT 0.73 0.35 1.06 1.01 ;
        RECT 2.575 1.3 2.915 1.63 ;
    END
    ANTENNADIFFAREA 0.5376 ;
    ANTENNAGATEAREA 0.279 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.018 LAYER li1 ;
  END QN

  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.35 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.279 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.088 LAYER li1 ;
  END S

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 1.23 0.085 1.56 0.84 ;
      RECT 2.28 0.085 2.705 0.5 ;
      RECT 0.23 0.085 0.56 0.84 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 1.115 2.29 1.445 3.245 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_udb_srlb_1
  
END LIBRARY
