# 
# LEF OUT 
# User Name : iptguser 
# Date : Mon Feb  4 15:39:15 2013
# 
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO scs8ls_macro_sync_posneg_nonret
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 15.36 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCD2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.645 4.51 12.08 5.135 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.144 LAYER li1 ;
  END SCD2

  PIN SCD1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.945 1.44 3.275 2.15 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14 LAYER li1 ;
  END SCD1

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.81 2.1 1.265 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.13 LAYER li1 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.075 3.68 1.405 6.31 ;
    END
    ANTENNADIFFAREA 0.5469 ;
    ANTENNAPARTIALMETALSIDEAREA 0.524 LAYER li1 ;
  END Q

  PIN SCO1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.91 1.82 15.27 2.98 ;
        RECT 15.1 1.13 15.27 1.82 ;
        RECT 14.915 0.35 15.27 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
    ANTENNAPARTIALMETALSIDEAREA 0.567 LAYER li1 ;
  END SCO1

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 15.36 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 15.36 6.905 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 15.36 3.575 ;
    END
  END vpwr

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 10.19 1.135 10.45 1.455 ;
        RECT 10.19 5.205 10.45 5.525 ;
        RECT 10.25 1.455 10.39 5.205 ;
    END
    PORT
      LAYER via ;
        RECT 10.245 1.22 10.395 1.37 ;
        RECT 10.245 5.29 10.395 5.44 ;
    END
    ANTENNAGATEAREA 0.558 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.101 LAYER met2 ;
  END CLK

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.79 1.875 8.05 2.195 ;
        RECT 7.79 4.835 8.05 5.155 ;
        RECT 7.85 2.195 7.99 4.835 ;
    END
    PORT
      LAYER via ;
        RECT 7.845 1.96 7.995 2.11 ;
        RECT 7.845 4.92 7.995 5.07 ;
    END
    ANTENNAGATEAREA 0.822 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.324 LAYER met2 ;
  END RESETB

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.59 1.505 12.85 1.825 ;
        RECT 12.59 5.205 12.85 5.525 ;
        RECT 12.65 1.825 12.79 5.205 ;
    END
    PORT
      LAYER via ;
        RECT 12.645 5.29 12.795 5.44 ;
        RECT 12.645 1.59 12.795 1.74 ;
    END
    ANTENNAGATEAREA 0.636 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.842 LAYER met2 ;
  END SCE

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 1.95 4.165 2.12 ;
      RECT 7.835 1.95 8.005 2.12 ;
      RECT 10.715 1.95 10.885 2.12 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 3.995 1.21 4.165 1.38 ;
      RECT 13.115 1.58 13.285 1.75 ;
      RECT 13.475 1.58 13.645 1.75 ;
      RECT 13.835 1.58 14.005 1.75 ;
      RECT 0.635 1.58 0.805 1.75 ;
      RECT 13.115 4.54 13.285 4.71 ;
      RECT 12.635 5.28 12.805 5.45 ;
      RECT 10.235 5.28 10.405 5.45 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 3.035 6.575 3.205 6.745 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 3.515 4.91 3.685 5.08 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 6.395 6.575 6.565 6.745 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 6.875 6.575 7.045 6.745 ;
      RECT 6.875 4.91 7.045 5.08 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 7.355 6.575 7.525 6.745 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.835 6.575 8.005 6.745 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 8.315 6.575 8.485 6.745 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 8.795 6.575 8.965 6.745 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 9.275 6.575 9.445 6.745 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 9.755 6.575 9.925 6.745 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 10.235 6.575 10.405 6.745 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 10.715 6.575 10.885 6.745 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 11.195 6.575 11.365 6.745 ;
      RECT 11.195 4.91 11.365 5.08 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 11.675 6.575 11.845 6.745 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 12.155 6.575 12.325 6.745 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 12.635 6.575 12.805 6.745 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 13.115 6.575 13.285 6.745 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 13.595 6.575 13.765 6.745 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 14.075 6.575 14.245 6.745 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 14.555 6.575 14.725 6.745 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 15.035 6.575 15.205 6.745 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
    LAYER via ;
      RECT 13.125 4.55 13.275 4.7 ;
      RECT 13.125 1.59 13.275 1.74 ;
    LAYER li1 ;
      RECT 6.71 1.03 6.88 2.32 ;
      RECT 7.495 1.26 8.315 1.575 ;
      RECT 6.14 0.86 6.88 1.03 ;
      RECT 6.14 0.595 6.47 0.86 ;
      RECT 8.725 1.715 9.005 2.755 ;
      RECT 8.725 1.09 8.895 1.715 ;
      RECT 7.05 0.92 8.895 1.09 ;
      RECT 7.05 1.09 7.325 1.805 ;
      RECT 8.27 0.595 8.655 0.92 ;
      RECT 10.145 1.955 10.315 2.55 ;
      RECT 9.585 1.785 10.315 1.955 ;
      RECT 9.29 2.55 10.315 2.88 ;
      RECT 9.585 1.265 9.755 1.785 ;
      RECT 9.585 1.095 11.395 1.265 ;
      RECT 9.585 0.77 9.755 1.095 ;
      RECT 11.065 1.265 11.395 1.275 ;
      RECT 9.405 0.35 9.755 0.77 ;
      RECT 9.985 1.445 11.735 1.615 ;
      RECT 9.985 1.435 10.315 1.445 ;
      RECT 11.14 1.615 11.31 2.52 ;
      RECT 11.565 0.925 11.735 1.445 ;
      RECT 10.945 2.52 11.31 2.98 ;
      RECT 11.01 0.755 11.735 0.925 ;
      RECT 11.01 0.35 11.34 0.755 ;
      RECT 7.835 1.815 8.165 2.15 ;
      RECT 10.64 1.82 10.97 2.15 ;
      RECT 14.57 1.3 14.93 1.63 ;
      RECT 13.91 2.12 14.24 2.98 ;
      RECT 13.91 1.95 14.74 2.12 ;
      RECT 14.57 1.63 14.74 1.95 ;
      RECT 14.57 1.28 14.74 1.3 ;
      RECT 13.555 1.11 14.74 1.28 ;
      RECT 13.555 0.8 14.235 1.11 ;
      RECT 12.995 0.35 13.325 1.13 ;
      RECT 13.565 1.75 14.35 1.78 ;
      RECT 13.565 1.45 14.35 1.58 ;
      RECT 13.07 1.58 14.35 1.75 ;
      RECT 13.07 1.75 13.325 2.98 ;
      RECT 13.07 1.13 13.325 1.58 ;
      RECT 11.98 2.1 12.31 2.98 ;
      RECT 12.085 1.63 12.31 2.1 ;
      RECT 12.085 1.3 12.87 1.63 ;
      RECT 12.085 0.35 12.335 1.3 ;
      RECT 2.085 3.68 2.44 4.975 ;
      RECT 2.07 4.975 2.44 5.305 ;
      RECT 2.085 5.305 2.44 6.31 ;
      RECT 5.315 4.52 6.19 4.69 ;
      RECT 5.315 3.68 6.085 4.52 ;
      RECT 6.02 4.69 6.19 5.36 ;
      RECT 5.87 5.36 7.735 5.53 ;
      RECT 7.405 4.79 7.735 5.36 ;
      RECT 2.985 4.54 4.025 4.71 ;
      RECT 2.985 4.71 3.315 5.62 ;
      RECT 3.855 4.71 4.025 4.78 ;
      RECT 2.985 5.62 4.885 5.79 ;
      RECT 3.855 4.78 5.145 4.95 ;
      RECT 4.715 5.79 4.885 6.04 ;
      RECT 4.815 3.68 5.145 4.78 ;
      RECT 4.715 6.04 5.69 6.37 ;
      RECT 2.645 4.37 2.815 5.96 ;
      RECT 2.645 4.2 4.445 4.37 ;
      RECT 2.645 5.96 3.19 6.21 ;
      RECT 4.195 4.37 4.445 4.61 ;
      RECT 3.17 3.68 3.5 4.2 ;
      RECT 6.36 4.52 6.975 4.69 ;
      RECT 6.805 4.385 6.975 4.52 ;
      RECT 6.36 4.69 6.655 5.19 ;
      RECT 6.805 4.215 8.425 4.385 ;
      RECT 7.95 4.385 8.12 5.565 ;
      RECT 6.805 3.68 7.135 4.215 ;
      RECT 8.095 3.68 8.425 4.215 ;
      RECT 7.95 5.565 8.215 5.895 ;
      RECT 9.865 4.525 10.445 4.84 ;
      RECT 9.865 4.84 10.035 5.04 ;
      RECT 9.705 5.04 10.035 5.37 ;
      RECT 9.865 5.37 10.035 5.62 ;
      RECT 9.865 5.62 10.635 5.79 ;
      RECT 11.2 3.86 13.475 4.03 ;
      RECT 10.805 5.475 12.16 5.645 ;
      RECT 12.66 3.7 13.475 3.86 ;
      RECT 11.99 5.645 12.16 5.895 ;
      RECT 11.99 5.895 12.925 6.065 ;
      RECT 8.625 4.185 11.45 4.355 ;
      RECT 8.625 3.68 8.875 4.185 ;
      RECT 10.805 4.355 11.45 4.36 ;
      RECT 11.2 4.03 11.45 4.185 ;
      RECT 10.805 4.36 10.975 5.475 ;
      RECT 11.2 3.68 11.45 3.86 ;
      RECT 10.805 5.645 10.975 5.96 ;
      RECT 8.725 5.96 10.975 6.13 ;
      RECT 8.725 5.565 8.975 5.96 ;
      RECT 8.29 4.555 9.535 4.84 ;
      RECT 9.105 4.525 9.535 4.555 ;
      RECT 8.29 4.84 8.62 4.885 ;
      RECT 9.205 4.84 9.535 5.225 ;
      RECT 8.385 5.225 9.535 5.395 ;
      RECT 8.385 5.395 8.555 6.115 ;
      RECT 9.205 5.395 9.535 5.79 ;
      RECT 7.61 6.115 8.555 6.405 ;
      RECT 7.61 5.87 7.78 6.115 ;
      RECT 5.055 5.7 7.78 5.87 ;
      RECT 5.055 5.46 5.385 5.7 ;
      RECT 12.335 4.37 12.665 5.08 ;
      RECT 12.335 4.2 14.765 4.37 ;
      RECT 14.515 4.37 14.765 5.42 ;
      RECT 14.515 3.68 14.765 4.2 ;
      RECT 13.26 5.42 14.765 5.61 ;
      RECT 13.26 5.61 13.59 5.725 ;
      RECT 14.435 5.61 14.765 6.24 ;
      RECT 12.9 4.54 13.795 4.88 ;
      RECT 14.015 4.58 14.345 5.08 ;
      RECT 12.835 5.08 14.345 5.25 ;
      RECT 12.33 5.25 13.005 5.705 ;
      RECT 4.485 5.29 4.815 5.435 ;
      RECT 4.485 5.19 5.7 5.29 ;
      RECT 4.485 5.12 5.85 5.19 ;
      RECT 5.53 4.86 5.85 5.12 ;
      RECT 3.485 5.12 3.885 5.45 ;
      RECT 3.485 4.88 3.685 5.12 ;
      RECT 10.205 5.11 10.605 5.45 ;
      RECT 6.845 4.86 7.195 5.19 ;
      RECT 11.145 4.635 11.475 5.305 ;
      RECT 11.49 6.235 13.715 6.405 ;
      RECT 13.385 5.895 13.715 6.235 ;
      RECT 11.49 5.815 11.82 6.235 ;
      RECT 0 3.245 15.36 3.415 ;
      RECT 14.41 2.29 14.74 3.245 ;
      RECT 11.48 2.1 11.81 3.245 ;
      RECT 12.54 1.82 12.87 3.245 ;
      RECT 11.735 3.415 12.065 3.69 ;
      RECT 13.985 3.415 14.315 4.03 ;
      RECT 8.385 1.745 8.555 3.245 ;
      RECT 2.67 3.415 3 4.03 ;
      RECT 3.67 3.415 4.275 4.01 ;
      RECT 4.705 2.73 5.035 3.245 ;
      RECT 3.095 2.685 3.425 3.245 ;
      RECT 6.255 3.415 6.585 4.35 ;
      RECT 7.335 3.415 7.585 4.045 ;
      RECT 9.555 3.415 9.885 4.015 ;
      RECT 7.205 2.66 7.54 3.245 ;
      RECT 10.485 2.52 10.735 3.245 ;
      RECT 10.64 3.415 10.97 4.015 ;
      RECT 1.575 3.415 1.905 4.84 ;
      RECT 0.615 2.345 0.945 3.245 ;
      RECT 1.575 5.53 1.905 6.575 ;
      RECT 3.68 5.98 4.15 6.575 ;
      RECT 9.715 6.3 10.075 6.575 ;
      RECT 6.66 6.04 6.99 6.575 ;
      RECT 10.815 6.3 11.305 6.575 ;
      RECT 13.935 5.78 14.265 6.575 ;
      RECT 0 6.575 15.36 6.745 ;
      RECT 0 -0.085 15.36 0.085 ;
      RECT 3.785 0.085 3.955 0.75 ;
      RECT 4.715 0.085 4.965 0.75 ;
      RECT 7.43 0.085 7.76 0.41 ;
      RECT 10.195 0.085 10.525 0.81 ;
      RECT 11.57 0.085 11.905 0.585 ;
      RECT 12.565 0.085 12.815 1.13 ;
      RECT 14.415 0.085 14.745 0.94 ;
      RECT 0.545 0.085 0.875 0.88 ;
      RECT 1.105 0.255 3.605 0.425 ;
      RECT 1.105 0.425 1.435 0.64 ;
      RECT 3.09 0.425 3.605 0.715 ;
      RECT 5.15 0.255 7.22 0.425 ;
      RECT 5.15 0.425 5.62 1.13 ;
      RECT 7.05 0.425 7.22 0.58 ;
      RECT 5.45 1.13 5.62 1.545 ;
      RECT 7.05 0.58 8.1 0.75 ;
      RECT 5.45 1.545 6.2 1.82 ;
      RECT 7.93 0.425 8.1 0.58 ;
      RECT 5.155 1.82 6.2 1.875 ;
      RECT 7.93 0.255 9.235 0.425 ;
      RECT 5.155 1.875 5.62 2.22 ;
      RECT 9.065 0.425 9.235 0.94 ;
      RECT 9.065 0.94 9.415 1.27 ;
      RECT 9.245 1.27 9.415 2.125 ;
      RECT 9.245 2.125 9.975 2.38 ;
      RECT 0.455 1.66 1.795 1.835 ;
      RECT 0.455 1.49 2.725 1.66 ;
      RECT 2.395 1.26 2.725 1.49 ;
      RECT 0.115 2.005 2.705 2.175 ;
      RECT 2.035 1.83 2.705 2.005 ;
      RECT 0.115 2.175 0.445 2.98 ;
      RECT 0.115 1.265 0.285 2.005 ;
      RECT 0.115 1.05 1.375 1.265 ;
      RECT 1.045 0.935 1.375 1.05 ;
      RECT 0.115 0.42 0.365 1.05 ;
      RECT 1.485 2.39 6.075 2.515 ;
      RECT 1.485 2.345 3.995 2.39 ;
      RECT 5.825 2.215 6.075 2.39 ;
      RECT 3.665 2.515 6.075 2.56 ;
      RECT 3.445 2.33 3.995 2.345 ;
      RECT 5.825 2.045 6.54 2.215 ;
      RECT 3.665 2.56 3.995 2.98 ;
      RECT 5.825 2.56 6.075 2.725 ;
      RECT 3.445 1.09 3.615 2.33 ;
      RECT 6.37 1.37 6.54 2.045 ;
      RECT 2.27 0.92 3.615 1.09 ;
      RECT 5.79 1.2 6.54 1.37 ;
      RECT 5.79 0.595 5.96 1.2 ;
      RECT 1.485 2.515 2.555 2.98 ;
      RECT 2.27 0.595 2.6 0.92 ;
      RECT 3.965 1.26 4.64 1.59 ;
      RECT 3.965 1.18 4.195 1.26 ;
      RECT 4.335 1.99 4.585 2.22 ;
      RECT 4.335 1.82 4.98 1.99 ;
      RECT 4.81 1.63 4.98 1.82 ;
      RECT 4.81 1.3 5.28 1.63 ;
      RECT 4.81 1.09 4.98 1.3 ;
      RECT 4.365 0.92 4.98 1.09 ;
      RECT 4.365 0.35 4.535 0.92 ;
      RECT 3.785 1.83 4.165 2.16 ;
      RECT 6.25 2.385 8.075 2.49 ;
      RECT 6.71 2.32 8.075 2.385 ;
      RECT 6.25 2.49 6.88 2.725 ;
      RECT 7.745 2.49 8.075 2.745 ;
      RECT 7.495 1.575 7.665 2.32 ;
    LAYER met2 ;
      RECT 13.07 1.505 13.33 1.825 ;
      RECT 13.13 1.665 13.27 4.625 ;
      RECT 13.07 4.465 13.33 4.785 ;
    LAYER met1 ;
      RECT 3.455 5.065 3.745 5.11 ;
      RECT 3.455 4.925 11.425 5.065 ;
      RECT 6.815 5.065 7.105 5.11 ;
      RECT 11.135 5.065 11.425 5.11 ;
      RECT 3.455 4.88 3.745 4.925 ;
      RECT 6.815 4.88 7.105 4.925 ;
      RECT 11.135 4.88 11.425 4.925 ;
      RECT 7.76 5.065 8.08 5.125 ;
      RECT 7.76 4.865 8.08 4.925 ;
      RECT 10.655 2.105 10.945 2.15 ;
      RECT 3.935 1.965 10.945 2.105 ;
      RECT 10.655 1.92 10.945 1.965 ;
      RECT 3.935 2.105 4.225 2.15 ;
      RECT 3.935 1.92 4.225 1.965 ;
      RECT 7.76 2.105 8.08 2.165 ;
      RECT 7.76 1.905 8.08 1.965 ;
      RECT 13.04 1.55 14.065 1.78 ;
      RECT 13.04 1.78 13.36 1.795 ;
      RECT 13.04 1.535 13.36 1.55 ;
      RECT 12.56 1.735 12.88 1.795 ;
      RECT 12.56 1.535 12.88 1.595 ;
      RECT 0.575 1.595 12.88 1.735 ;
      RECT 0.575 1.735 0.865 1.78 ;
      RECT 0.575 1.55 0.865 1.595 ;
      RECT 10.16 1.365 10.48 1.425 ;
      RECT 10.16 1.165 10.48 1.225 ;
      RECT 3.935 1.225 10.48 1.365 ;
      RECT 3.935 1.365 4.225 1.41 ;
      RECT 3.935 1.18 4.225 1.225 ;
      RECT 13.04 4.495 13.36 4.755 ;
      RECT 12.56 5.235 12.88 5.495 ;
      RECT 10.16 5.235 10.48 5.495 ;
  END
END scs8ls_macro_sync_posneg_nonret

MACRO scs8ls_macro_sync_posneg_ret
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 20.64 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCD2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.85 4.54 16.195 5.055 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.104 LAYER li1 ;
  END SCD2

  PIN SCD1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.35 1.55 3.715 1.88 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.071 LAYER li1 ;
  END SCD1

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.84 2.135 2.17 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.112 LAYER li1 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585 3.585 0.925 6.395 ;
    END
    ANTENNADIFFAREA 0.5301 ;
    ANTENNAPARTIALMETALSIDEAREA 0.562 LAYER li1 ;
  END Q

  PIN SCO1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.81 5.53 19.165 6.31 ;
        RECT 18.81 4.84 18.98 5.53 ;
        RECT 18.81 3.68 19.17 4.84 ;
    END
    ANTENNADIFFAREA 0.5413 ;
    ANTENNAPARTIALMETALSIDEAREA 0.567 LAYER li1 ;
  END SCO1

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 20.57 2.945 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 3.715 20.57 3.985 ;
        RECT 10.175 3.985 10.465 4 ;
        RECT 10.655 3.985 10.945 4 ;
    END
    PORT
      LAYER via ;
        RECT 10.245 2.74 10.395 2.89 ;
        RECT 11.685 2.74 11.835 2.89 ;
        RECT 11.685 3.77 11.835 3.92 ;
        RECT 10.245 3.77 10.395 3.92 ;
    END
  END kapwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 20.64 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 20.64 6.905 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 20.64 3.575 ;
    END
  END vpwr

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.67 1.505 10.93 1.825 ;
        RECT 10.67 5.205 10.93 5.525 ;
        RECT 10.73 1.825 10.87 5.205 ;
    END
    PORT
      LAYER via ;
        RECT 10.725 5.29 10.875 5.44 ;
        RECT 10.725 1.59 10.875 1.74 ;
    END
    ANTENNAGATEAREA 1.196 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.842 LAYER met2 ;
  END RESETB

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.35 1.135 18.61 1.455 ;
        RECT 18.35 5.575 18.61 5.895 ;
        RECT 18.41 1.455 18.55 5.575 ;
    END
    PORT
      LAYER via ;
        RECT 18.405 5.66 18.555 5.81 ;
        RECT 18.405 1.22 18.555 1.37 ;
    END
    ANTENNAGATEAREA 1.196 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.36 LAYER met2 ;
  END SLEEPB

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 11.15 4.82 11.41 5.14 ;
        RECT 11.15 1.505 11.41 1.825 ;
        RECT 11.21 1.825 11.35 4.82 ;
    END
    PORT
      LAYER via ;
        RECT 11.205 4.905 11.355 5.055 ;
        RECT 11.205 1.59 11.355 1.74 ;
    END
    ANTENNAGATEAREA 0.318 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5725 LAYER met2 ;
  END CLK

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.99 1.135 15.25 1.455 ;
        RECT 14.99 5.205 15.25 5.525 ;
        RECT 15.05 1.455 15.19 5.205 ;
    END
    PORT
      LAYER via ;
        RECT 15.045 5.29 15.195 5.44 ;
        RECT 15.045 1.22 15.195 1.37 ;
    END
    ANTENNAGATEAREA 0.636 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.101 LAYER met2 ;
  END SCE

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 15.515 6.575 15.685 6.745 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.995 6.575 16.165 6.745 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 16.475 6.575 16.645 6.745 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 16.955 6.575 17.125 6.745 ;
      RECT 16.955 3.245 17.125 3.415 ;
      RECT 17.435 6.575 17.605 6.745 ;
      RECT 17.435 3.245 17.605 3.415 ;
      RECT 17.915 6.575 18.085 6.745 ;
      RECT 17.915 3.245 18.085 3.415 ;
      RECT 18.395 6.575 18.565 6.745 ;
      RECT 18.395 3.245 18.565 3.415 ;
      RECT 6.875 3.775 7.045 3.945 ;
      RECT 18.875 6.575 19.045 6.745 ;
      RECT 19.355 6.575 19.525 6.745 ;
      RECT 19.835 6.575 20.005 6.745 ;
      RECT 20.315 6.575 20.485 6.745 ;
      RECT 18.875 3.245 19.045 3.415 ;
      RECT 19.355 3.245 19.525 3.415 ;
      RECT 19.835 3.245 20.005 3.415 ;
      RECT 20.315 3.245 20.485 3.415 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 7.355 4.91 7.525 5.08 ;
      RECT 8.315 4.91 8.485 5.08 ;
      RECT 11.54 5.28 11.71 5.45 ;
      RECT 16.955 4.91 17.125 5.08 ;
      RECT 17.915 5.28 18.085 5.45 ;
      RECT 20.315 4.91 20.485 5.08 ;
      RECT 20.315 1.95 20.485 2.12 ;
      RECT 18.38 1.21 18.55 1.38 ;
      RECT 16.955 1.58 17.125 1.75 ;
      RECT 0.635 1.58 0.805 1.75 ;
      RECT 3.995 1.58 4.165 1.75 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 15.035 2.735 15.205 2.905 ;
      RECT 15.515 2.735 15.685 2.905 ;
      RECT 17.435 2.735 17.605 2.905 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.835 6.575 8.005 6.745 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 8.315 6.575 8.485 6.745 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 8.795 6.575 8.965 6.745 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 9.275 6.575 9.445 6.745 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 9.755 6.575 9.925 6.745 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 10.235 6.575 10.405 6.745 ;
      RECT 10.235 3.8 10.405 3.97 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 6.875 6.575 7.045 6.745 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 3.035 6.575 3.205 6.745 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 6.395 6.575 6.565 6.745 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 4.475 4.54 4.645 4.71 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 7.355 6.575 7.525 6.745 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 10.715 6.575 10.885 6.745 ;
      RECT 10.715 3.8 10.885 3.97 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 11.195 6.575 11.365 6.745 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 11.675 6.575 11.845 6.745 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 12.155 6.575 12.325 6.745 ;
      RECT 12.155 4.54 12.325 4.71 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 12.635 6.575 12.805 6.745 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 13.115 6.575 13.285 6.745 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 13.595 6.575 13.765 6.745 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 14.075 6.575 14.245 6.745 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 14.555 6.575 14.725 6.745 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 15.035 6.575 15.205 6.745 ;
      RECT 15.035 4.54 15.205 4.71 ;
      RECT 15.995 2.735 16.165 2.905 ;
      RECT 20.315 -0.085 20.485 0.085 ;
      RECT 20.315 3.245 20.485 3.415 ;
      RECT 19.835 -0.085 20.005 0.085 ;
      RECT 19.835 3.245 20.005 3.415 ;
      RECT 19.355 -0.085 19.525 0.085 ;
      RECT 19.355 3.245 19.525 3.415 ;
      RECT 18.875 -0.085 19.045 0.085 ;
      RECT 18.875 3.245 19.045 3.415 ;
      RECT 18.395 -0.085 18.565 0.085 ;
      RECT 18.395 3.245 18.565 3.415 ;
      RECT 17.915 -0.085 18.085 0.085 ;
      RECT 17.915 3.245 18.085 3.415 ;
      RECT 17.435 -0.085 17.605 0.085 ;
      RECT 17.435 3.245 17.605 3.415 ;
      RECT 16.955 -0.085 17.125 0.085 ;
      RECT 16.955 2.735 17.125 2.905 ;
      RECT 16.955 3.245 17.125 3.415 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 16.475 2.735 16.645 2.905 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 2.735 14.725 2.905 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
    LAYER li1 ;
      RECT 8.705 5.275 10.025 5.445 ;
      RECT 9.695 5.16 10.025 5.275 ;
      RECT 6.64 4.65 7.525 4.71 ;
      RECT 6.64 4.54 8.215 4.65 ;
      RECT 6.64 4.71 6.81 5.115 ;
      RECT 7.695 4.65 7.865 5.395 ;
      RECT 7.255 4.48 8.215 4.54 ;
      RECT 5.575 5.115 6.81 5.285 ;
      RECT 7.695 5.395 8.3 5.645 ;
      RECT 8.045 3.935 8.215 4.48 ;
      RECT 7.255 3.925 7.525 4.48 ;
      RECT 5.575 4.925 5.97 5.115 ;
      RECT 8.045 3.765 9.31 3.935 ;
      RECT 9.14 3.935 9.31 4.14 ;
      RECT 9.14 4.14 11.645 4.31 ;
      RECT 11.475 3.755 11.645 4.14 ;
      RECT 11.475 3.585 13.51 3.755 ;
      RECT 13.34 3.755 13.51 4.725 ;
      RECT 13.34 4.725 13.67 5.055 ;
      RECT 6.67 3.755 7.075 4.37 ;
      RECT 6.67 3.585 7.875 3.755 ;
      RECT 7.705 3.755 7.875 4.31 ;
      RECT 8.385 4.48 11.985 4.65 ;
      RECT 8.385 4.105 8.64 4.48 ;
      RECT 10.535 4.65 11.985 4.71 ;
      RECT 11.815 4.34 11.985 4.48 ;
      RECT 11.815 4.17 13.065 4.34 ;
      RECT 12.735 4.34 13.065 5.26 ;
      RECT 12.735 3.925 13.065 4.17 ;
      RECT 12.735 5.26 13.205 5.51 ;
      RECT 9.48 3.64 10.435 3.97 ;
      RECT 10.685 3.585 11.305 3.97 ;
      RECT 15.46 4.2 17.1 4.37 ;
      RECT 16.77 3.585 17.1 4.2 ;
      RECT 15.51 5.225 16.66 5.395 ;
      RECT 16.49 5.395 16.66 5.735 ;
      RECT 16.49 5.735 17.22 6.065 ;
      RECT 13.915 4.555 14.085 4.755 ;
      RECT 13.755 3.905 14.085 4.555 ;
      RECT 13.915 4.755 14.775 4.925 ;
      RECT 14.605 3.755 14.775 4.755 ;
      RECT 13.915 4.925 14.085 5.225 ;
      RECT 14.605 3.585 15.63 3.755 ;
      RECT 13.375 5.225 14.085 5.395 ;
      RECT 15.46 3.755 15.63 4.2 ;
      RECT 13.375 5.395 13.545 5.68 ;
      RECT 12.05 5.68 13.545 5.85 ;
      RECT 15.51 4.37 15.68 5.225 ;
      RECT 12.05 5.28 12.38 5.68 ;
      RECT 12.155 4.51 12.565 5.11 ;
      RECT 14.985 3.925 15.235 5.065 ;
      RECT 14.985 5.065 15.34 5.395 ;
      RECT 16.41 4.54 18.615 4.71 ;
      RECT 18.11 3.585 18.615 4.54 ;
      RECT 16.41 4.71 16.745 4.75 ;
      RECT 18.365 4.71 18.615 6.375 ;
      RECT 19.34 4.54 20.17 4.71 ;
      RECT 19.84 3.68 20.17 4.54 ;
      RECT 19.34 4.71 19.51 5.03 ;
      RECT 19.15 5.03 19.51 5.36 ;
      RECT 19.34 5.36 19.51 5.38 ;
      RECT 19.34 5.38 20.525 5.55 ;
      RECT 19.845 5.55 20.525 5.86 ;
      RECT 9.86 6.125 10.145 6.315 ;
      RECT 9.86 5.955 11.165 6.125 ;
      RECT 10.835 6.125 11.165 6.295 ;
      RECT 7.16 4.88 7.525 5.365 ;
      RECT 8.035 4.82 8.515 5.105 ;
      RECT 11.54 6.235 14.115 6.405 ;
      RECT 11.54 5.05 11.71 6.235 ;
      RECT 10.58 4.88 11.71 5.05 ;
      RECT 10.58 5.05 10.98 5.445 ;
      RECT 14.02 5.735 14.35 6.065 ;
      RECT 14.02 5.565 16.32 5.735 ;
      RECT 16.15 5.735 16.32 6.065 ;
      RECT 16.915 4.88 17.635 5.48 ;
      RECT 17.805 4.88 18.135 5.565 ;
      RECT 15.64 6.235 17.65 6.405 ;
      RECT 15.64 5.905 15.97 6.235 ;
      RECT 17.4 5.735 17.65 6.235 ;
      RECT 19.73 4.88 20.515 5.21 ;
      RECT 5.035 0.595 6.055 0.765 ;
      RECT 5.035 0.765 5.205 1.25 ;
      RECT 5.725 0.765 6.055 1.265 ;
      RECT 4.545 1.25 5.205 1.42 ;
      RECT 4.545 1.42 4.715 2.07 ;
      RECT 2.98 2.07 4.715 2.1 ;
      RECT 2.305 2.1 4.755 2.24 ;
      RECT 4.47 2.24 4.755 2.99 ;
      RECT 2.305 2.24 3.08 2.325 ;
      RECT 2.305 2.325 2.635 2.34 ;
      RECT 1.225 2.34 2.635 2.51 ;
      RECT 1.96 2.51 2.635 2.99 ;
      RECT 1.225 1.5 2.08 1.67 ;
      RECT 1.83 0.935 2.08 1.5 ;
      RECT 1.225 1.67 1.395 2.34 ;
      RECT 14.985 0.425 15.315 0.6 ;
      RECT 14.985 0.255 17.1 0.425 ;
      RECT 14.015 0.6 15.315 0.77 ;
      RECT 16.93 0.425 17.1 0.78 ;
      RECT 14.015 0.77 14.185 1.32 ;
      RECT 16.93 0.78 18.345 0.95 ;
      RECT 12.93 1.32 14.185 1.5 ;
      RECT 18.015 0.345 18.345 0.78 ;
      RECT 17.895 0.95 18.065 1.85 ;
      RECT 17.895 1.85 18.49 2.18 ;
      RECT 11.905 0.575 12.235 1.155 ;
      RECT 11.1 1.155 12.235 1.325 ;
      RECT 11.1 1.325 11.43 2.01 ;
      RECT 11.1 2.01 16.08 2.18 ;
      RECT 14.695 1.93 16.08 2.01 ;
      RECT 14.695 1.28 14.955 1.93 ;
      RECT 12.695 0.575 12.945 0.98 ;
      RECT 12.695 0.98 13.845 1.15 ;
      RECT 13.675 0.575 13.845 0.98 ;
      RECT 20.205 0.35 20.535 1.82 ;
      RECT 19.995 1.82 20.535 2.155 ;
      RECT 19.995 2.155 20.325 2.975 ;
      RECT 19.235 0.345 19.685 0.975 ;
      RECT 18.735 0.975 19.685 1.145 ;
      RECT 18.735 1.145 18.905 1.815 ;
      RECT 19.515 1.145 19.685 1.315 ;
      RECT 18.735 1.815 18.985 2.18 ;
      RECT 19.515 1.315 20.02 1.645 ;
      RECT 16.105 0.595 16.435 0.94 ;
      RECT 14.355 0.94 16.435 0.95 ;
      RECT 14.355 0.95 16.76 1.11 ;
      RECT 14.355 1.11 14.525 1.67 ;
      RECT 16.105 1.11 16.76 1.12 ;
      RECT 11.64 1.67 14.525 1.84 ;
      RECT 16.59 1.12 17.495 1.29 ;
      RECT 11.64 1.51 11.97 1.67 ;
      RECT 17.325 1.29 17.495 2.01 ;
      RECT 16.855 2.01 17.495 2.18 ;
      RECT 3.92 1.55 4.25 1.88 ;
      RECT 0.605 1.5 0.935 2.17 ;
      RECT 4.925 1.92 5.095 2.6 ;
      RECT 4.885 1.59 5.215 1.92 ;
      RECT 4.925 2.6 5.95 2.77 ;
      RECT 5.78 2.435 7.68 2.6 ;
      RECT 5.78 2.43 8.725 2.435 ;
      RECT 8.395 2.435 8.725 2.825 ;
      RECT 7.51 2.265 8.725 2.43 ;
      RECT 8.555 2.825 8.725 2.905 ;
      RECT 8.395 1.665 8.725 2.265 ;
      RECT 8.555 2.905 13.455 3.075 ;
      RECT 8.395 1.495 9.4 1.665 ;
      RECT 13.125 2.745 13.455 2.905 ;
      RECT 9.07 1.665 9.4 1.825 ;
      RECT 8.395 1.335 8.99 1.495 ;
      RECT 5.265 2.26 5.555 2.43 ;
      RECT 5.265 2.09 7.11 2.26 ;
      RECT 6.78 1.675 7.11 2.09 ;
      RECT 5.385 1.265 5.555 2.09 ;
      RECT 6.78 1.345 7.795 1.675 ;
      RECT 5.375 0.935 5.555 1.265 ;
      RECT 14.525 2.69 17.73 3.025 ;
      RECT 18.235 1.12 18.565 1.45 ;
      RECT 16.59 1.46 17.155 1.79 ;
      RECT 3.41 3.755 3.74 4.135 ;
      RECT 3.41 3.585 5.97 3.755 ;
      RECT 5.64 3.755 5.97 4.415 ;
      RECT 4.135 4.655 4.305 4.865 ;
      RECT 4.02 4.865 4.305 5.035 ;
      RECT 4.02 5.035 4.19 6.235 ;
      RECT 4.02 6.235 6.295 6.405 ;
      RECT 5.065 6.08 5.395 6.235 ;
      RECT 6.125 6.045 6.295 6.235 ;
      RECT 6.125 5.875 7.185 6.045 ;
      RECT 7.015 6.045 7.185 6.155 ;
      RECT 7.015 6.155 9.215 6.325 ;
      RECT 9.045 5.785 9.215 6.155 ;
      RECT 9.045 5.615 11.37 5.785 ;
      RECT 10.195 4.99 10.365 5.615 ;
      RECT 11.15 5.22 11.37 5.615 ;
      RECT 8.76 4.82 10.365 4.99 ;
      RECT 8.76 4.99 9.09 5.07 ;
      RECT 4.475 4.51 4.645 5.205 ;
      RECT 4.36 5.205 4.645 5.535 ;
      RECT 1.55 4.225 1.74 5.015 ;
      RECT 1.55 3.585 1.88 4.225 ;
      RECT 1.095 5.015 1.74 5.345 ;
      RECT 1.57 5.345 1.74 5.935 ;
      RECT 1.57 5.935 1.9 6.265 ;
      RECT 3.68 4.475 3.85 5.385 ;
      RECT 3.68 4.34 4.08 4.475 ;
      RECT 2.93 5.385 3.85 5.555 ;
      RECT 3.68 4.305 5.065 4.34 ;
      RECT 2.93 5.555 3.1 6.235 ;
      RECT 4.815 4.34 5.065 5.705 ;
      RECT 3.91 4.165 5.065 4.305 ;
      RECT 2.07 6.235 3.1 6.405 ;
      RECT 4.565 5.705 5.065 5.875 ;
      RECT 2.07 5.765 2.24 6.235 ;
      RECT 4.565 5.875 4.895 6.065 ;
      RECT 1.91 5.095 2.24 5.765 ;
      RECT 2.515 4.525 3.51 4.855 ;
      RECT 2.515 3.905 2.835 4.525 ;
      RECT 2.515 4.855 2.685 5.725 ;
      RECT 2.415 5.725 2.685 6.065 ;
      RECT 5.235 4.585 6.47 4.755 ;
      RECT 5.235 4.755 5.405 5.535 ;
      RECT 6.14 4.755 6.47 4.945 ;
      RECT 5.235 5.535 7.525 5.705 ;
      RECT 5.625 5.705 5.955 6.065 ;
      RECT 7.355 5.705 7.525 5.815 ;
      RECT 7.355 5.815 8.875 5.985 ;
      RECT 8.705 5.445 8.875 5.815 ;
      RECT 0 -0.085 20.64 0.085 ;
      RECT 0.535 0.085 0.865 0.99 ;
      RECT 3.615 0.085 3.865 1.04 ;
      RECT 7.05 0.085 7.38 0.835 ;
      RECT 8.02 0.085 8.35 0.825 ;
      RECT 11.365 0.085 11.695 0.985 ;
      RECT 13.125 0.085 13.455 0.81 ;
      RECT 17.475 0.085 17.805 0.61 ;
      RECT 18.805 0.085 19.055 0.805 ;
      RECT 19.855 0.085 20.025 1.13 ;
      RECT 0 3.245 20.64 3.415 ;
      RECT 19.495 1.815 19.825 3.245 ;
      RECT 19.34 3.415 19.67 4.37 ;
      RECT 15.8 3.415 16.05 4.03 ;
      RECT 17.61 3.415 17.94 4.225 ;
      RECT 3.245 2.41 4.3 3.245 ;
      RECT 7.85 2.605 8.18 3.245 ;
      RECT 6.12 2.77 6.45 3.245 ;
      RECT 14.265 3.415 14.435 4.585 ;
      RECT 2.085 3.415 2.335 4.365 ;
      RECT 3.005 3.415 3.24 4.355 ;
      RECT 0.645 2.34 0.975 3.245 ;
      RECT 1.095 3.415 1.345 4.34 ;
      RECT 12.21 2.35 19.325 2.52 ;
      RECT 12.21 2.52 12.54 2.565 ;
      RECT 13.625 2.52 13.955 2.97 ;
      RECT 16.25 1.74 16.42 2.35 ;
      RECT 19.155 1.645 19.325 2.35 ;
      RECT 9.835 2.565 12.54 2.735 ;
      RECT 15.985 1.41 16.42 1.74 ;
      RECT 19.075 1.315 19.345 1.645 ;
      RECT 9.835 2.04 10.5 2.565 ;
      RECT 10.19 0.605 10.5 2.04 ;
      RECT 19.335 5.72 19.665 6.575 ;
      RECT 0 6.575 20.64 6.745 ;
      RECT 3.27 5.725 3.6 6.575 ;
      RECT 1.105 5.515 1.355 6.575 ;
      RECT 6.56 6.215 6.81 6.575 ;
      RECT 9.385 6 9.69 6.575 ;
      RECT 10.315 6.295 10.645 6.575 ;
      RECT 14.555 5.905 14.885 6.575 ;
      RECT 17.855 5.945 18.185 6.575 ;
      RECT 1.07 0.425 1.32 0.99 ;
      RECT 1.07 0.255 3.405 0.425 ;
      RECT 3.155 0.425 3.405 1.04 ;
      RECT 4.615 0.425 4.865 1.08 ;
      RECT 4.615 0.255 6.59 0.425 ;
      RECT 6.26 0.425 6.59 0.835 ;
      RECT 4.045 0.58 4.375 1.21 ;
      RECT 2.645 1.21 4.375 1.38 ;
      RECT 2.645 0.74 2.975 1.21 ;
      RECT 1.49 0.595 2.475 0.765 ;
      RECT 2.305 0.765 2.475 1.6 ;
      RECT 1.49 0.765 1.66 1.16 ;
      RECT 2.305 1.6 2.88 1.93 ;
      RECT 0.105 1.16 1.66 1.33 ;
      RECT 0.105 0.53 0.355 1.16 ;
      RECT 0.105 1.33 0.435 2.99 ;
      RECT 9.2 0.435 9.53 0.995 ;
      RECT 9.2 0.265 10.93 0.435 ;
      RECT 7.59 0.995 9.53 1.005 ;
      RECT 10.68 0.435 10.93 2.395 ;
      RECT 7.59 0.575 7.84 0.995 ;
      RECT 6.28 1.005 9.53 1.165 ;
      RECT 6.28 1.165 8.135 1.175 ;
      RECT 9.2 1.165 9.53 1.285 ;
      RECT 6.28 1.175 6.61 1.485 ;
      RECT 7.965 1.175 8.135 1.845 ;
      RECT 7.32 1.845 8.135 2.095 ;
    LAYER via ;
      RECT 20.325 4.92 20.475 5.07 ;
      RECT 20.325 1.96 20.475 2.11 ;
    LAYER met2 ;
      RECT 10.19 3.685 10.45 4.005 ;
      RECT 10.19 2.655 10.45 2.975 ;
      RECT 10.25 2.975 10.39 3.685 ;
      RECT 11.63 2.655 11.89 2.975 ;
      RECT 11.63 3.685 11.89 4.005 ;
      RECT 11.69 2.975 11.83 3.685 ;
      RECT 20.27 4.835 20.53 5.155 ;
      RECT 20.27 1.875 20.53 2.195 ;
      RECT 20.33 2.195 20.47 4.835 ;
    LAYER met1 ;
      RECT 4.415 4.695 4.705 4.74 ;
      RECT 4.415 4.555 15.265 4.695 ;
      RECT 12.095 4.695 12.385 4.74 ;
      RECT 14.975 4.695 15.265 4.74 ;
      RECT 4.415 4.51 4.705 4.555 ;
      RECT 12.095 4.51 12.385 4.555 ;
      RECT 14.975 4.51 15.265 4.555 ;
      RECT 18.32 1.165 18.64 1.425 ;
      RECT 0.575 1.55 0.865 1.78 ;
      RECT 0.65 1.225 15.28 1.365 ;
      RECT 14.96 1.365 15.28 1.425 ;
      RECT 14.96 1.165 15.28 1.225 ;
      RECT 0.65 1.365 0.79 1.55 ;
      RECT 8.255 5.065 8.545 5.11 ;
      RECT 8.255 4.88 8.545 4.925 ;
      RECT 8.255 4.925 11.44 5.065 ;
      RECT 11.12 5.065 11.44 5.11 ;
      RECT 11.12 4.85 11.44 4.925 ;
      RECT 7.295 4.88 7.585 5.11 ;
      RECT 7.37 5.11 7.51 5.665 ;
      RECT 18.32 5.805 18.64 5.865 ;
      RECT 7.37 5.665 18.64 5.805 ;
      RECT 18.32 5.605 18.64 5.665 ;
      RECT 11.48 5.435 11.77 5.48 ;
      RECT 11.48 5.25 11.77 5.295 ;
      RECT 10.64 5.295 11.77 5.435 ;
      RECT 10.64 5.435 10.96 5.495 ;
      RECT 10.64 5.235 10.96 5.295 ;
      RECT 16.895 1.735 17.185 1.78 ;
      RECT 16.895 1.55 17.185 1.595 ;
      RECT 11.12 1.595 17.185 1.735 ;
      RECT 11.12 1.735 11.44 1.795 ;
      RECT 11.12 1.535 11.44 1.595 ;
      RECT 3.935 1.735 4.225 1.78 ;
      RECT 3.935 1.55 4.225 1.595 ;
      RECT 3.935 1.595 10.96 1.735 ;
      RECT 10.64 1.735 10.96 1.795 ;
      RECT 10.64 1.535 10.96 1.595 ;
      RECT 17.855 5.435 18.145 5.48 ;
      RECT 17.855 5.25 18.145 5.295 ;
      RECT 14.96 5.295 18.145 5.435 ;
      RECT 14.96 5.435 15.28 5.495 ;
      RECT 14.96 5.235 15.28 5.295 ;
      RECT 16.895 5.065 17.185 5.11 ;
      RECT 16.895 4.88 17.185 4.925 ;
      RECT 16.895 4.925 20.56 5.065 ;
      RECT 20.24 5.065 20.56 5.125 ;
      RECT 20.24 4.865 20.56 4.925 ;
      RECT 20.24 1.905 20.56 2.165 ;
  END
END scs8ls_macro_sync_posneg_ret

MACRO scs8ls_macro_sync_pospos_nonret
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 14.88 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455 1.66 1.795 1.835 ;
        RECT 0.455 1.49 2.725 1.66 ;
        RECT 2.395 1.26 2.725 1.49 ;
    END
    ANTENNAGATEAREA 0.318 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.501 LAYER li1 ;
  END SCE

  PIN SCD1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.945 1.44 3.275 2.15 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14 LAYER li1 ;
  END SCD1

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.81 2.1 1.265 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.13 LAYER li1 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 3.68 0.37 5.53 ;
        RECT 0.115 5.53 0.445 6.31 ;
    END
    ANTENNADIFFAREA 0.5413 ;
    ANTENNAPARTIALMETALSIDEAREA 0.524 LAYER li1 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.88 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 14.88 6.905 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.88 3.575 ;
    END
  END vpwr

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 9.23 1.135 9.49 1.455 ;
        RECT 9.23 5.205 9.49 5.525 ;
        RECT 9.29 1.455 9.43 5.205 ;
    END
    PORT
      LAYER via ;
        RECT 9.285 5.29 9.435 5.44 ;
        RECT 9.285 1.22 9.435 1.37 ;
    END
    ANTENNAGATEAREA 0.558 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.101 LAYER met2 ;
  END CLK

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.79 1.875 8.05 2.195 ;
        RECT 7.79 4.465 8.05 4.785 ;
        RECT 7.85 2.195 7.99 4.465 ;
    END
    PORT
      LAYER via ;
        RECT 7.845 4.55 7.995 4.7 ;
        RECT 7.845 1.96 7.995 2.11 ;
    END
    ANTENNAGATEAREA 0.822 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.065 LAYER met2 ;
  END RESETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 7.835 1.95 8.005 2.12 ;
      RECT 10.715 1.95 10.885 2.12 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 13.115 1.95 13.285 2.12 ;
      RECT 13.595 4.91 13.765 5.08 ;
      RECT 12.155 4.91 12.325 5.08 ;
      RECT 11.675 5.65 11.845 5.82 ;
      RECT 10.235 4.91 10.405 5.08 ;
      RECT 9.275 5.28 9.445 5.45 ;
      RECT 3.995 1.21 4.165 1.38 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 3.035 6.575 3.205 6.745 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 6.395 6.575 6.565 6.745 ;
      RECT 6.875 6.575 7.045 6.745 ;
      RECT 7.355 6.575 7.525 6.745 ;
      RECT 7.835 6.575 8.005 6.745 ;
      RECT 8.315 6.575 8.485 6.745 ;
      RECT 8.795 6.575 8.965 6.745 ;
      RECT 9.275 6.575 9.445 6.745 ;
      RECT 9.755 6.575 9.925 6.745 ;
      RECT 10.235 6.575 10.405 6.745 ;
      RECT 10.715 6.575 10.885 6.745 ;
      RECT 11.195 6.575 11.365 6.745 ;
      RECT 11.675 6.575 11.845 6.745 ;
      RECT 12.155 6.575 12.325 6.745 ;
      RECT 12.635 6.575 12.805 6.745 ;
      RECT 13.115 6.575 13.285 6.745 ;
      RECT 9.275 4.54 9.445 4.71 ;
      RECT 5.435 4.54 5.605 4.71 ;
      RECT 2.555 4.54 2.725 4.71 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 13.595 6.575 13.765 6.745 ;
      RECT 14.075 6.575 14.245 6.745 ;
      RECT 14.555 6.575 14.725 6.745 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 1.95 4.165 2.12 ;
    LAYER li1 ;
      RECT 5.15 0.255 7.22 0.425 ;
      RECT 7.05 0.425 7.22 0.58 ;
      RECT 7.05 0.58 8.1 0.75 ;
      RECT 7.93 0.425 8.1 0.58 ;
      RECT 7.93 0.255 9.235 0.425 ;
      RECT 9.065 0.425 9.235 0.94 ;
      RECT 9.065 0.94 9.415 1.27 ;
      RECT 9.245 1.27 9.415 2.125 ;
      RECT 9.245 2.125 9.975 2.38 ;
      RECT 3.785 1.83 4.165 2.16 ;
      RECT 6.14 0.86 6.88 1.03 ;
      RECT 6.14 0.595 6.47 0.86 ;
      RECT 6.71 1.03 6.88 2.32 ;
      RECT 6.71 2.32 8.075 2.385 ;
      RECT 7.495 1.575 7.665 2.32 ;
      RECT 6.25 2.385 8.075 2.49 ;
      RECT 7.495 1.26 8.315 1.575 ;
      RECT 6.25 2.49 6.88 2.725 ;
      RECT 7.745 2.49 8.075 2.745 ;
      RECT 8.725 1.715 9.005 2.755 ;
      RECT 8.725 1.09 8.895 1.715 ;
      RECT 7.05 0.92 8.895 1.09 ;
      RECT 7.05 1.09 7.325 1.805 ;
      RECT 8.27 0.595 8.655 0.92 ;
      RECT 10.145 1.955 10.315 2.55 ;
      RECT 9.585 1.785 10.315 1.955 ;
      RECT 9.29 2.55 10.315 2.88 ;
      RECT 9.585 1.265 9.755 1.785 ;
      RECT 9.585 1.095 11.395 1.265 ;
      RECT 9.585 0.77 9.755 1.095 ;
      RECT 11.065 1.265 11.395 1.275 ;
      RECT 9.405 0.35 9.755 0.77 ;
      RECT 9.985 1.445 11.735 1.615 ;
      RECT 9.985 1.435 10.315 1.445 ;
      RECT 11.14 1.615 11.31 2.52 ;
      RECT 11.565 0.925 11.735 1.445 ;
      RECT 10.945 2.52 11.31 2.98 ;
      RECT 11.01 0.755 11.735 0.925 ;
      RECT 11.01 0.35 11.34 0.755 ;
      RECT 7.835 1.815 8.165 2.15 ;
      RECT 13.07 1.13 13.325 2.98 ;
      RECT 12.995 0.35 13.325 1.13 ;
      RECT 11.98 2.1 12.31 2.98 ;
      RECT 12.085 1.63 12.31 2.1 ;
      RECT 12.085 1.3 12.87 1.63 ;
      RECT 12.085 0.35 12.335 1.3 ;
      RECT 10.64 1.82 10.97 2.15 ;
      RECT 1.13 3.68 1.46 4.56 ;
      RECT 1.13 4.56 1.355 5.03 ;
      RECT 0.57 5.03 1.355 5.36 ;
      RECT 1.105 5.36 1.355 6.31 ;
      RECT 4.435 3.905 4.715 4.945 ;
      RECT 4.545 4.945 4.715 5.57 ;
      RECT 4.545 5.57 6.39 5.74 ;
      RECT 4.785 5.74 5.17 6.065 ;
      RECT 6.115 4.855 6.39 5.57 ;
      RECT 3.125 4.11 3.295 4.705 ;
      RECT 3.125 3.78 4.15 4.11 ;
      RECT 3.125 4.705 3.855 4.875 ;
      RECT 3.685 4.875 3.855 5.395 ;
      RECT 2.045 5.395 3.855 5.565 ;
      RECT 3.685 5.565 3.855 5.89 ;
      RECT 2.045 5.385 2.375 5.395 ;
      RECT 3.685 5.89 4.035 6.31 ;
      RECT 3.465 4.28 4.195 4.535 ;
      RECT 4.025 4.535 4.195 5.39 ;
      RECT 4.025 5.39 4.375 5.72 ;
      RECT 4.205 5.72 4.375 6.235 ;
      RECT 4.205 6.235 5.51 6.405 ;
      RECT 5.34 6.08 5.51 6.235 ;
      RECT 5.34 5.91 6.39 6.08 ;
      RECT 6.22 6.08 6.39 6.235 ;
      RECT 6.22 6.235 8.29 6.405 ;
      RECT 7.82 5.53 8.29 6.235 ;
      RECT 7.82 5.115 7.99 5.53 ;
      RECT 7.24 4.84 7.99 5.115 ;
      RECT 7.24 4.785 8.285 4.84 ;
      RECT 7.82 4.44 8.285 4.785 ;
      RECT 5.775 4.34 5.945 5.085 ;
      RECT 5.365 4.275 6.73 4.34 ;
      RECT 5.125 5.085 5.945 5.4 ;
      RECT 5.365 4.17 7.19 4.275 ;
      RECT 6.56 4.34 6.73 5.63 ;
      RECT 5.365 3.915 5.695 4.17 ;
      RECT 6.56 3.935 7.19 4.17 ;
      RECT 6.56 5.63 7.3 5.8 ;
      RECT 6.97 5.8 7.3 6.065 ;
      RECT 2.13 4.14 2.3 5.045 ;
      RECT 2.13 3.68 2.495 4.14 ;
      RECT 1.705 5.045 3.455 5.215 ;
      RECT 1.705 5.215 1.875 5.735 ;
      RECT 3.125 5.215 3.455 5.225 ;
      RECT 1.705 5.735 2.43 5.905 ;
      RECT 2.1 5.905 2.43 6.31 ;
      RECT 8.855 4.44 9.105 4.67 ;
      RECT 8.46 4.67 9.105 4.84 ;
      RECT 8.46 4.84 8.63 5.03 ;
      RECT 8.16 5.03 8.63 5.36 ;
      RECT 8.46 5.36 8.63 5.57 ;
      RECT 8.46 5.57 9.075 5.74 ;
      RECT 8.905 5.74 9.075 6.31 ;
      RECT 9.275 4.5 9.655 4.83 ;
      RECT 10.735 4.485 13.325 4.655 ;
      RECT 12.995 3.68 13.325 4.485 ;
      RECT 10.735 4.655 11.405 4.83 ;
      RECT 13.155 4.655 13.325 5.395 ;
      RECT 12.065 5.395 13.325 5.61 ;
      RECT 12.065 5.61 12.395 5.725 ;
      RECT 13.075 5.61 13.325 6.24 ;
      RECT 13.525 4.175 13.825 5.665 ;
      RECT 13.525 3.585 14.055 4.175 ;
      RECT 14.485 4.325 14.795 5.815 ;
      RECT 14.265 5.815 14.795 6.405 ;
      RECT 5.275 4.51 5.605 4.845 ;
      RECT 2.47 4.51 2.8 4.84 ;
      RECT 10.165 4.51 10.495 5.22 ;
      RECT 9.245 5.4 9.475 5.48 ;
      RECT 8.8 5.07 9.475 5.4 ;
      RECT 9.835 6.235 12.335 6.405 ;
      RECT 9.835 5.945 10.35 6.235 ;
      RECT 12.005 6.02 12.335 6.235 ;
      RECT 11.34 5.395 11.875 5.85 ;
      RECT 10.715 5 12.985 5.17 ;
      RECT 11.645 4.825 12.985 5 ;
      RECT 10.715 5.17 11.045 5.4 ;
      RECT 7.365 4.145 11.955 4.27 ;
      RECT 7.365 4.27 7.615 4.445 ;
      RECT 9.445 4.27 11.955 4.315 ;
      RECT 7.365 4.1 9.775 4.145 ;
      RECT 10.885 3.68 11.955 4.145 ;
      RECT 6.9 4.445 7.615 4.615 ;
      RECT 9.445 4.315 9.995 4.33 ;
      RECT 7.365 3.935 7.615 4.1 ;
      RECT 9.445 3.68 9.775 4.1 ;
      RECT 6.9 4.615 7.07 5.29 ;
      RECT 9.825 4.33 9.995 5.57 ;
      RECT 6.9 5.29 7.65 5.46 ;
      RECT 9.825 5.57 11.17 5.74 ;
      RECT 7.48 5.46 7.65 6.065 ;
      RECT 10.84 5.74 11.17 6.065 ;
      RECT 8.385 1.745 8.555 3.245 ;
      RECT 11.48 2.1 11.81 3.245 ;
      RECT 12.54 1.82 12.87 3.245 ;
      RECT 2.705 3.415 2.955 4.14 ;
      RECT 4.885 3.415 5.055 4.915 ;
      RECT 5.9 3.415 6.235 4 ;
      RECT 4.705 2.73 5.035 3.245 ;
      RECT 3.095 2.685 3.425 3.245 ;
      RECT 8.405 3.415 8.735 3.93 ;
      RECT 10.015 3.415 10.345 3.975 ;
      RECT 7.205 2.66 7.54 3.245 ;
      RECT 10.485 2.52 10.735 3.245 ;
      RECT 12.495 3.415 12.825 4.315 ;
      RECT 14.265 3.415 14.595 4.155 ;
      RECT 0 3.245 14.88 3.415 ;
      RECT 0.57 3.415 0.9 4.84 ;
      RECT 0.615 2.345 0.945 3.245 ;
      RECT 1.63 3.415 1.96 4.56 ;
      RECT 1.535 6.075 1.87 6.575 ;
      RECT 0.625 5.53 0.875 6.575 ;
      RECT 5.68 6.25 6.01 6.575 ;
      RECT 2.915 5.85 3.245 6.575 ;
      RECT 8.475 5.91 8.725 6.575 ;
      RECT 9.485 5.91 9.655 6.575 ;
      RECT 12.565 5.78 12.895 6.575 ;
      RECT 13.725 5.835 14.055 6.575 ;
      RECT 0 6.575 14.88 6.745 ;
      RECT 1.485 2.39 6.075 2.515 ;
      RECT 5.825 2.215 6.075 2.39 ;
      RECT 1.485 2.345 3.995 2.39 ;
      RECT 3.665 2.515 6.075 2.56 ;
      RECT 5.825 2.045 6.54 2.215 ;
      RECT 3.445 2.33 3.995 2.345 ;
      RECT 3.665 2.56 3.995 2.98 ;
      RECT 5.825 2.56 6.075 2.725 ;
      RECT 6.37 1.37 6.54 2.045 ;
      RECT 3.445 1.09 3.615 2.33 ;
      RECT 5.79 1.2 6.54 1.37 ;
      RECT 2.27 0.92 3.615 1.09 ;
      RECT 5.79 0.595 5.96 1.2 ;
      RECT 1.485 2.515 2.555 2.98 ;
      RECT 2.27 0.595 2.6 0.92 ;
      RECT 3.785 0.085 3.955 0.75 ;
      RECT 4.715 0.085 4.965 0.75 ;
      RECT 7.43 0.085 7.76 0.41 ;
      RECT 10.195 0.085 10.525 0.81 ;
      RECT 11.57 0.085 11.905 0.585 ;
      RECT 12.565 0.085 12.815 1.13 ;
      RECT 0 -0.085 14.88 0.085 ;
      RECT 0.545 0.085 0.875 0.88 ;
      RECT 1.105 0.425 1.435 0.64 ;
      RECT 1.105 0.255 3.605 0.425 ;
      RECT 3.09 0.425 3.605 0.715 ;
      RECT 0.115 2.005 2.705 2.175 ;
      RECT 2.035 1.83 2.705 2.005 ;
      RECT 0.115 2.175 0.445 2.98 ;
      RECT 0.115 1.265 0.285 2.005 ;
      RECT 0.115 0.42 0.365 1.05 ;
      RECT 0.115 1.05 1.375 1.265 ;
      RECT 1.045 0.935 1.375 1.05 ;
      RECT 3.965 1.26 4.64 1.59 ;
      RECT 3.965 1.18 4.195 1.26 ;
      RECT 4.335 1.99 4.585 2.22 ;
      RECT 4.335 1.82 4.98 1.99 ;
      RECT 4.81 1.63 4.98 1.82 ;
      RECT 4.81 1.3 5.28 1.63 ;
      RECT 4.81 1.09 4.98 1.3 ;
      RECT 4.365 0.92 4.98 1.09 ;
      RECT 4.365 0.35 4.535 0.92 ;
      RECT 5.155 1.875 5.62 2.22 ;
      RECT 5.155 1.82 6.2 1.875 ;
      RECT 5.45 1.545 6.2 1.82 ;
      RECT 5.45 1.13 5.62 1.545 ;
      RECT 5.15 0.425 5.62 1.13 ;
    LAYER via ;
      RECT 11.685 1.96 11.835 2.11 ;
      RECT 11.685 5.66 11.835 5.81 ;
    LAYER met2 ;
      RECT 11.63 1.875 11.89 2.195 ;
      RECT 11.69 2.035 11.83 5.735 ;
      RECT 11.63 5.575 11.89 5.895 ;
    LAYER met1 ;
      RECT 2.495 4.695 2.785 4.74 ;
      RECT 2.495 4.555 9.505 4.695 ;
      RECT 2.495 4.51 2.785 4.555 ;
      RECT 5.375 4.695 5.665 4.74 ;
      RECT 9.215 4.695 9.505 4.74 ;
      RECT 5.375 4.51 5.665 4.555 ;
      RECT 9.215 4.51 9.505 4.555 ;
      RECT 7.76 4.695 8.08 4.755 ;
      RECT 7.76 4.495 8.08 4.555 ;
      RECT 10.655 2.105 10.945 2.15 ;
      RECT 3.935 1.965 10.945 2.105 ;
      RECT 10.655 1.92 10.945 1.965 ;
      RECT 3.935 2.105 4.225 2.15 ;
      RECT 3.935 1.92 4.225 1.965 ;
      RECT 7.76 2.105 8.08 2.165 ;
      RECT 7.76 1.905 8.08 1.965 ;
      RECT 11.6 2.105 11.92 2.165 ;
      RECT 11.6 1.905 11.92 1.965 ;
      RECT 11.6 1.965 13.345 2.105 ;
      RECT 13.055 2.105 13.345 2.15 ;
      RECT 13.055 1.92 13.345 1.965 ;
      RECT 11.6 5.605 11.92 5.865 ;
      RECT 9.2 5.235 9.52 5.495 ;
      RECT 9.2 1.365 9.52 1.425 ;
      RECT 9.2 1.165 9.52 1.225 ;
      RECT 3.935 1.225 9.52 1.365 ;
      RECT 3.935 1.365 4.225 1.41 ;
      RECT 3.935 1.18 4.225 1.225 ;
      RECT 10.175 5.065 10.465 5.11 ;
      RECT 10.175 4.88 10.465 4.925 ;
      RECT 10.175 4.925 13.825 5.065 ;
      RECT 13.535 5.065 13.825 5.11 ;
      RECT 13.535 4.88 13.825 4.925 ;
      RECT 12.095 5.065 12.385 5.11 ;
      RECT 12.095 4.88 12.385 4.925 ;
  END
END scs8ls_macro_sync_pospos_nonret

MACRO scs8ls_macro_sync_pospos_ret
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 22.08 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCD1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.35 1.55 3.715 1.88 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.071 LAYER li1 ;
  END SCD1

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.84 2.135 2.17 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.112 LAYER li1 ;
  END D

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 4.84 0.435 6.31 ;
        RECT 0.105 4.505 0.645 4.84 ;
        RECT 0.315 3.685 0.645 4.505 ;
    END
    ANTENNADIFFAREA 0.5395 ;
    ANTENNAPARTIALMETALSIDEAREA 0.565 LAYER li1 ;
  END Q

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.5 0.935 2.17 ;
    END
    ANTENNAGATEAREA 0.318 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.132 LAYER li1 ;
  END SCE

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 22.01 2.945 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 3.715 22.01 3.985 ;
    END
    PORT
      LAYER via ;
        RECT 10.245 3.77 10.395 3.92 ;
        RECT 11.685 3.77 11.835 3.92 ;
        RECT 11.685 2.74 11.835 2.89 ;
        RECT 10.245 2.74 10.395 2.89 ;
    END
  END kapwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 22.08 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 22.08 6.905 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 22.08 3.575 ;
    END
  END vpwr

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.67 1.505 10.93 1.825 ;
        RECT 10.67 5.205 10.93 5.525 ;
        RECT 10.73 1.825 10.87 5.205 ;
    END
    PORT
      LAYER via ;
        RECT 10.725 1.59 10.875 1.74 ;
        RECT 10.725 5.29 10.875 5.44 ;
    END
    ANTENNAGATEAREA 1.196 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.842 LAYER met2 ;
  END RESETB

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.35 1.135 18.61 1.455 ;
        RECT 18.35 5.575 18.61 5.895 ;
        RECT 18.41 1.455 18.55 5.575 ;
    END
    PORT
      LAYER via ;
        RECT 18.405 1.22 18.555 1.37 ;
        RECT 18.405 5.66 18.555 5.81 ;
    END
    ANTENNAGATEAREA 1.196 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.36 LAYER met2 ;
  END SLEEPB

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 11.15 4.82 11.41 5.14 ;
        RECT 11.15 1.505 11.41 1.825 ;
        RECT 11.21 1.825 11.35 4.82 ;
    END
    PORT
      LAYER via ;
        RECT 11.205 1.59 11.355 1.74 ;
        RECT 11.205 4.905 11.355 5.055 ;
    END
    ANTENNAGATEAREA 0.318 LAYER met2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5725 LAYER met2 ;
  END CLK

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 16.955 3.245 17.125 3.415 ;
      RECT 17.435 6.575 17.605 6.745 ;
      RECT 17.435 3.245 17.605 3.415 ;
      RECT 20.795 6.575 20.965 6.745 ;
      RECT 21.275 6.575 21.445 6.745 ;
      RECT 21.755 6.575 21.925 6.745 ;
      RECT 20.795 3.245 20.965 3.415 ;
      RECT 21.275 3.245 21.445 3.415 ;
      RECT 21.755 3.245 21.925 3.415 ;
      RECT 20.795 -0.085 20.965 0.085 ;
      RECT 20.795 3.245 20.965 3.415 ;
      RECT 21.755 3.245 21.925 3.415 ;
      RECT 21.755 -0.085 21.925 0.085 ;
      RECT 21.275 -0.085 21.445 0.085 ;
      RECT 21.275 3.245 21.445 3.415 ;
      RECT 16.955 1.58 17.125 1.75 ;
      RECT 18.38 1.21 18.55 1.38 ;
      RECT 20.315 1.95 20.485 2.12 ;
      RECT 20.795 4.91 20.965 5.08 ;
      RECT 19.835 4.91 20.005 5.08 ;
      RECT 18.875 4.54 19.045 4.71 ;
      RECT 16.955 4.91 17.125 5.08 ;
      RECT 16.475 4.91 16.645 5.08 ;
      RECT 2.075 5.28 2.245 5.45 ;
      RECT 3.515 4.91 3.685 5.08 ;
      RECT 3.995 1.58 4.165 1.75 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 15.035 2.735 15.205 2.905 ;
      RECT 15.515 2.735 15.685 2.905 ;
      RECT 17.435 2.735 17.605 2.905 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 3.035 6.575 3.205 6.745 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 3.515 3.755 3.685 3.925 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 3.995 3.755 4.165 3.925 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 5.915 3.755 6.085 3.925 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 6.395 6.575 6.565 6.745 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 6.875 6.575 7.045 6.745 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 7.355 6.575 7.525 6.745 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.835 6.575 8.005 6.745 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 8.315 6.575 8.485 6.745 ;
      RECT 17.915 6.575 18.085 6.745 ;
      RECT 17.915 3.245 18.085 3.415 ;
      RECT 18.395 6.575 18.565 6.745 ;
      RECT 18.395 3.245 18.565 3.415 ;
      RECT 18.875 6.575 19.045 6.745 ;
      RECT 18.875 3.245 19.045 3.415 ;
      RECT 19.355 6.575 19.525 6.745 ;
      RECT 19.355 3.245 19.525 3.415 ;
      RECT 19.835 6.575 20.005 6.745 ;
      RECT 19.835 3.245 20.005 3.415 ;
      RECT 20.315 6.575 20.485 6.745 ;
      RECT 20.315 3.245 20.485 3.415 ;
      RECT 5.435 3.755 5.605 3.925 ;
      RECT 4.955 3.755 5.125 3.925 ;
      RECT 3.035 3.755 3.205 3.925 ;
      RECT 4.475 3.755 4.645 3.925 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 8.795 6.575 8.965 6.745 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 9.275 6.575 9.445 6.745 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 9.755 6.575 9.925 6.745 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 10.235 6.575 10.405 6.745 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 10.715 6.575 10.885 6.745 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 11.195 6.575 11.365 6.745 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 11.675 6.575 11.845 6.745 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 12.155 6.575 12.325 6.745 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 12.635 6.575 12.805 6.745 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 13.115 6.575 13.285 6.745 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 13.595 6.575 13.765 6.745 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 14.075 6.575 14.245 6.745 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 14.555 6.575 14.725 6.745 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 15.035 6.575 15.205 6.745 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 15.515 6.575 15.685 6.745 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.995 6.575 16.165 6.745 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 16.475 6.575 16.645 6.745 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 16.955 6.575 17.125 6.745 ;
      RECT 15.995 2.735 16.165 2.905 ;
      RECT 20.315 -0.085 20.485 0.085 ;
      RECT 20.315 3.245 20.485 3.415 ;
      RECT 19.835 -0.085 20.005 0.085 ;
      RECT 19.835 3.245 20.005 3.415 ;
      RECT 19.355 -0.085 19.525 0.085 ;
      RECT 19.355 3.245 19.525 3.415 ;
      RECT 18.875 -0.085 19.045 0.085 ;
      RECT 18.875 3.245 19.045 3.415 ;
      RECT 18.395 -0.085 18.565 0.085 ;
      RECT 18.395 3.245 18.565 3.415 ;
      RECT 17.915 -0.085 18.085 0.085 ;
      RECT 17.915 3.245 18.085 3.415 ;
      RECT 17.435 -0.085 17.605 0.085 ;
      RECT 17.435 3.245 17.605 3.415 ;
      RECT 16.955 -0.085 17.125 0.085 ;
      RECT 16.955 2.735 17.125 2.905 ;
      RECT 16.955 3.245 17.125 3.415 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 16.475 2.735 16.645 2.905 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 2.735 14.725 2.905 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
    LAYER li1 ;
      RECT 11.11 5.655 13.05 5.665 ;
      RECT 11.11 5.495 14.36 5.655 ;
      RECT 12.8 5.665 13.05 6.085 ;
      RECT 11.11 5.375 11.44 5.495 ;
      RECT 12.505 5.485 14.36 5.495 ;
      RECT 14.03 5.175 14.36 5.485 ;
      RECT 12.505 4.815 12.675 5.485 ;
      RECT 12.505 4.565 13.32 4.815 ;
      RECT 14.525 2.69 17.73 3.025 ;
      RECT 13.53 4.57 13.86 4.985 ;
      RECT 13.53 4.4 15.375 4.57 ;
      RECT 12.845 4.985 13.86 5.315 ;
      RECT 15.085 4.57 15.255 5.395 ;
      RECT 15.085 4.23 15.375 4.4 ;
      RECT 15.085 5.395 15.265 5.725 ;
      RECT 15.925 4.59 16.095 5.24 ;
      RECT 15.925 4.56 17.66 4.59 ;
      RECT 15.435 5.24 16.095 5.41 ;
      RECT 15.885 4.42 18.335 4.56 ;
      RECT 15.435 5.41 15.605 5.895 ;
      RECT 15.885 3.67 16.17 4.42 ;
      RECT 17.56 4.335 18.335 4.42 ;
      RECT 14.585 5.895 15.605 6.065 ;
      RECT 18.005 4.32 18.335 4.335 ;
      RECT 14.585 5.395 14.915 5.895 ;
      RECT 18.005 4.15 19.415 4.32 ;
      RECT 19.245 4.32 19.415 4.99 ;
      RECT 18.005 3.67 18.68 4.15 ;
      RECT 18.56 4.99 19.415 5.16 ;
      RECT 18.56 5.16 18.81 5.725 ;
      RECT 20.205 3.67 20.535 5.33 ;
      RECT 18.98 5.33 20.535 5.5 ;
      RECT 18.98 5.5 19.15 5.895 ;
      RECT 20.285 5.5 20.535 6.13 ;
      RECT 18.165 5.895 19.15 6.065 ;
      RECT 18.165 5.06 18.335 5.895 ;
      RECT 17.76 4.73 18.335 5.06 ;
      RECT 18.505 4.49 19.075 4.82 ;
      RECT 19.705 4.49 20.035 5.16 ;
      RECT 21.685 4.325 21.995 5.815 ;
      RECT 21.465 5.815 21.995 6.405 ;
      RECT 20.725 3.585 21.255 4.175 ;
      RECT 20.725 4.175 21.025 5.665 ;
      RECT 2.075 5.21 2.405 5.54 ;
      RECT 3.485 4.87 4.05 5.2 ;
      RECT 6.795 5.68 6.965 6.085 ;
      RECT 6.795 5.51 7.945 5.68 ;
      RECT 7.695 5.68 7.945 6.085 ;
      RECT 14.05 6.235 16.025 6.405 ;
      RECT 14.05 5.825 14.38 6.235 ;
      RECT 15.775 5.58 16.025 6.235 ;
      RECT 16.265 5.45 16.595 6.08 ;
      RECT 16.265 5.28 17.995 5.45 ;
      RECT 17.665 5.45 17.995 5.92 ;
      RECT 16.39 4.78 16.72 5.11 ;
      RECT 16.925 4.78 17.29 5.11 ;
      RECT 17.235 6.235 19.57 6.405 ;
      RECT 19.32 5.67 19.57 6.235 ;
      RECT 17.235 5.62 17.485 6.235 ;
      RECT 14.015 0.6 15.315 0.77 ;
      RECT 16.93 0.425 17.1 0.78 ;
      RECT 14.015 0.77 14.185 1.32 ;
      RECT 16.93 0.78 18.345 0.95 ;
      RECT 12.93 1.32 14.185 1.5 ;
      RECT 18.015 0.345 18.345 0.78 ;
      RECT 17.895 0.95 18.065 1.85 ;
      RECT 17.895 1.85 18.49 2.18 ;
      RECT 20.205 0.35 20.535 1.82 ;
      RECT 19.995 1.82 20.535 2.155 ;
      RECT 19.995 2.155 20.325 2.975 ;
      RECT 19.235 0.345 19.685 0.975 ;
      RECT 18.735 0.975 19.685 1.145 ;
      RECT 18.735 1.145 18.905 1.815 ;
      RECT 19.515 1.145 19.685 1.315 ;
      RECT 18.735 1.815 18.985 2.18 ;
      RECT 19.515 1.315 20.02 1.645 ;
      RECT 4.045 0.58 4.375 1.21 ;
      RECT 2.645 1.21 4.375 1.38 ;
      RECT 2.645 0.74 2.975 1.21 ;
      RECT 4.925 2.6 5.95 2.77 ;
      RECT 4.925 1.92 5.095 2.6 ;
      RECT 5.78 2.435 7.68 2.6 ;
      RECT 4.885 1.59 5.215 1.92 ;
      RECT 5.78 2.43 8.725 2.435 ;
      RECT 8.395 2.435 8.725 2.825 ;
      RECT 7.51 2.265 8.725 2.43 ;
      RECT 8.555 2.825 8.725 2.905 ;
      RECT 8.395 1.665 8.725 2.265 ;
      RECT 8.555 2.905 13.455 3.075 ;
      RECT 8.395 1.495 9.4 1.665 ;
      RECT 13.125 2.745 13.455 2.905 ;
      RECT 9.07 1.665 9.4 1.825 ;
      RECT 8.395 1.335 8.99 1.495 ;
      RECT 2.305 2.1 4.755 2.24 ;
      RECT 4.47 2.24 4.755 2.99 ;
      RECT 2.98 2.07 4.715 2.1 ;
      RECT 4.545 1.42 4.715 2.07 ;
      RECT 4.545 1.25 5.205 1.42 ;
      RECT 5.035 0.765 5.205 1.25 ;
      RECT 5.035 0.595 6.055 0.765 ;
      RECT 5.725 0.765 6.055 1.265 ;
      RECT 1.96 2.51 2.635 2.99 ;
      RECT 1.225 2.34 2.635 2.51 ;
      RECT 2.305 2.325 2.635 2.34 ;
      RECT 2.305 2.24 3.08 2.325 ;
      RECT 1.225 1.5 2.08 1.67 ;
      RECT 1.83 0.935 2.08 1.5 ;
      RECT 1.225 1.67 1.395 2.34 ;
      RECT 3.92 1.55 4.25 1.88 ;
      RECT 5.265 2.26 5.555 2.43 ;
      RECT 5.265 2.09 7.11 2.26 ;
      RECT 5.385 1.265 5.555 2.09 ;
      RECT 6.78 1.675 7.11 2.09 ;
      RECT 5.375 0.935 5.555 1.265 ;
      RECT 6.78 1.345 7.795 1.675 ;
      RECT 11.905 0.575 12.235 1.155 ;
      RECT 11.1 1.155 12.235 1.325 ;
      RECT 11.1 1.325 11.43 2.01 ;
      RECT 11.1 2.01 16.08 2.18 ;
      RECT 14.695 1.93 16.08 2.01 ;
      RECT 14.695 1.28 14.955 1.93 ;
      RECT 12.695 0.575 12.945 0.98 ;
      RECT 12.695 0.98 13.845 1.15 ;
      RECT 13.675 0.575 13.845 0.98 ;
      RECT 11.64 1.67 14.525 1.84 ;
      RECT 11.64 1.51 11.97 1.67 ;
      RECT 14.355 1.11 14.525 1.67 ;
      RECT 14.355 0.95 16.76 1.11 ;
      RECT 16.105 1.11 16.76 1.12 ;
      RECT 14.355 0.94 16.435 0.95 ;
      RECT 16.59 1.12 17.495 1.29 ;
      RECT 16.105 0.595 16.435 0.94 ;
      RECT 17.325 1.29 17.495 2.01 ;
      RECT 16.855 2.01 17.495 2.18 ;
      RECT 16.59 1.46 17.155 1.79 ;
      RECT 18.235 1.12 18.565 1.45 ;
      RECT 1.655 4.48 1.905 4.845 ;
      RECT 1.735 4.845 1.905 5.515 ;
      RECT 0.955 5.515 1.905 5.685 ;
      RECT 0.955 5.685 1.405 6.315 ;
      RECT 0.955 5.345 1.125 5.515 ;
      RECT 0.62 5.015 1.125 5.345 ;
      RECT 2.15 4.48 2.745 4.81 ;
      RECT 2.575 4.81 2.745 5.71 ;
      RECT 2.295 5.71 3.71 5.88 ;
      RECT 2.295 5.88 2.625 6.315 ;
      RECT 3.54 5.88 3.71 6.235 ;
      RECT 3.54 6.235 5.655 6.405 ;
      RECT 5.325 6.06 5.655 6.235 ;
      RECT 5.325 5.89 6.625 6.06 ;
      RECT 6.455 5.34 6.625 5.89 ;
      RECT 6.455 5.16 7.71 5.34 ;
      RECT 3.145 4.65 3.315 5.37 ;
      RECT 3.145 4.48 3.785 4.65 ;
      RECT 3.145 5.37 4.05 5.54 ;
      RECT 3.88 5.54 4.535 5.55 ;
      RECT 3.88 5.55 6.285 5.71 ;
      RECT 4.205 5.71 6.285 5.72 ;
      RECT 6.115 4.99 6.285 5.55 ;
      RECT 4.205 5.72 4.535 6.065 ;
      RECT 6.115 4.82 9 4.99 ;
      RECT 8.67 4.99 9 5.15 ;
      RECT 4.56 4.65 5.945 4.73 ;
      RECT 4.56 4.48 9.54 4.65 ;
      RECT 5.685 4.73 5.945 5.38 ;
      RECT 9.21 4.65 9.54 5.335 ;
      RECT 8.405 5.335 9.54 5.505 ;
      RECT 8.405 5.505 8.735 6.085 ;
      RECT 2.91 3.635 6.115 3.97 ;
      RECT 7.185 3.755 7.515 3.915 ;
      RECT 7.185 3.585 12.085 3.755 ;
      RECT 11.915 3.755 12.085 3.835 ;
      RECT 11.915 3.835 12.245 4.225 ;
      RECT 11.915 4.225 14.86 4.23 ;
      RECT 11.915 4.23 13.13 4.395 ;
      RECT 12.96 4.06 14.86 4.225 ;
      RECT 11.915 4.395 12.245 4.995 ;
      RECT 14.69 3.89 15.715 4.06 ;
      RECT 11.24 4.995 12.245 5.165 ;
      RECT 15.545 4.06 15.715 4.74 ;
      RECT 11.65 5.165 12.245 5.325 ;
      RECT 11.24 4.835 11.57 4.995 ;
      RECT 15.425 4.74 15.755 5.07 ;
      RECT 9.71 4.265 9.96 6.225 ;
      RECT 9.71 6.225 11.44 6.395 ;
      RECT 11.11 5.665 11.44 6.225 ;
      RECT 0.535 0.085 0.865 0.99 ;
      RECT 3.615 0.085 3.865 1.04 ;
      RECT 7.05 0.085 7.38 0.835 ;
      RECT 8.02 0.085 8.35 0.825 ;
      RECT 11.365 0.085 11.695 0.985 ;
      RECT 13.125 0.085 13.455 0.81 ;
      RECT 17.475 0.085 17.805 0.61 ;
      RECT 18.805 0.085 19.055 0.805 ;
      RECT 19.855 0.085 20.025 1.13 ;
      RECT 0 -0.085 22.08 0.085 ;
      RECT 3.245 2.41 4.3 3.245 ;
      RECT 7.85 2.605 8.18 3.245 ;
      RECT 19.495 1.815 19.825 3.245 ;
      RECT 6.12 2.77 6.45 3.245 ;
      RECT 12.46 3.415 12.79 4.055 ;
      RECT 14.19 3.415 14.52 3.89 ;
      RECT 16.34 3.415 17.395 4.25 ;
      RECT 19.665 3.415 19.995 4.32 ;
      RECT 21.465 3.415 21.795 4.155 ;
      RECT 0 3.245 22.08 3.415 ;
      RECT 0.645 2.34 0.975 3.245 ;
      RECT 0.815 3.415 1.145 4.845 ;
      RECT 12.21 2.35 19.325 2.52 ;
      RECT 12.21 2.52 12.54 2.565 ;
      RECT 13.625 2.52 13.955 2.97 ;
      RECT 16.25 1.74 16.42 2.35 ;
      RECT 19.155 1.645 19.325 2.35 ;
      RECT 9.835 2.565 12.54 2.735 ;
      RECT 15.985 1.41 16.42 1.74 ;
      RECT 19.075 1.315 19.345 1.645 ;
      RECT 9.835 2.04 10.5 2.565 ;
      RECT 10.19 0.605 10.5 2.04 ;
      RECT 2.835 6.05 3.165 6.575 ;
      RECT 1.585 5.855 1.835 6.575 ;
      RECT 0.615 5.53 0.785 6.575 ;
      RECT 7.185 5.85 7.515 6.575 ;
      RECT 8.945 5.675 9.275 6.575 ;
      RECT 12.29 5.835 12.62 6.575 ;
      RECT 13.26 5.825 13.59 6.575 ;
      RECT 19.775 5.67 20.105 6.575 ;
      RECT 16.775 5.62 17.025 6.575 ;
      RECT 20.925 5.835 21.255 6.575 ;
      RECT 0 6.575 22.08 6.745 ;
      RECT 1.315 4.14 8.43 4.31 ;
      RECT 1.315 4.31 1.485 5.015 ;
      RECT 4.22 4.31 4.39 4.92 ;
      RECT 8.1 4.095 8.43 4.14 ;
      RECT 6.685 3.69 7.015 4.14 ;
      RECT 1.295 5.015 1.565 5.345 ;
      RECT 4.22 4.92 4.655 5.25 ;
      RECT 8.1 3.925 10.805 4.095 ;
      RECT 10.14 4.095 10.805 4.62 ;
      RECT 10.14 4.62 10.45 6.055 ;
      RECT 0.105 1.16 1.66 1.33 ;
      RECT 1.49 0.765 1.66 1.16 ;
      RECT 1.49 0.595 2.475 0.765 ;
      RECT 2.305 0.765 2.475 1.6 ;
      RECT 2.305 1.6 2.88 1.93 ;
      RECT 0.105 0.53 0.355 1.16 ;
      RECT 0.105 1.33 0.435 2.99 ;
      RECT 4.615 0.425 4.865 1.08 ;
      RECT 4.615 0.255 6.59 0.425 ;
      RECT 6.26 0.425 6.59 0.835 ;
      RECT 1.07 0.425 1.32 0.99 ;
      RECT 1.07 0.255 3.405 0.425 ;
      RECT 3.155 0.425 3.405 1.04 ;
      RECT 9.2 0.435 9.53 0.995 ;
      RECT 9.2 0.265 10.93 0.435 ;
      RECT 7.59 0.995 9.53 1.005 ;
      RECT 10.68 0.435 10.93 2.395 ;
      RECT 7.59 0.575 7.84 0.995 ;
      RECT 6.28 1.005 9.53 1.165 ;
      RECT 6.28 1.165 8.135 1.175 ;
      RECT 9.2 1.165 9.53 1.285 ;
      RECT 6.28 1.175 6.61 1.485 ;
      RECT 7.965 1.175 8.135 1.845 ;
      RECT 7.32 1.845 8.135 2.095 ;
      RECT 14.985 0.425 15.315 0.6 ;
      RECT 14.985 0.255 17.1 0.425 ;
    LAYER via ;
      RECT 20.325 1.96 20.475 2.11 ;
      RECT 20.325 4.55 20.475 4.7 ;
    LAYER met2 ;
      RECT 10.19 3.685 10.45 4.005 ;
      RECT 10.19 2.655 10.45 2.975 ;
      RECT 10.25 2.975 10.39 3.685 ;
      RECT 11.63 2.655 11.89 2.975 ;
      RECT 11.63 3.685 11.89 4.005 ;
      RECT 11.69 2.975 11.83 3.685 ;
      RECT 20.27 1.875 20.53 2.195 ;
      RECT 20.27 4.465 20.53 4.785 ;
      RECT 20.33 2.195 20.47 4.465 ;
    LAYER met1 ;
      RECT 18.815 4.695 19.105 4.74 ;
      RECT 18.815 4.51 19.105 4.555 ;
      RECT 18.815 4.555 20.56 4.695 ;
      RECT 20.24 4.695 20.56 4.755 ;
      RECT 20.24 4.495 20.56 4.555 ;
      RECT 19.775 5.065 20.065 5.11 ;
      RECT 19.775 4.88 20.065 4.925 ;
      RECT 16.895 5.065 17.185 5.11 ;
      RECT 16.895 4.88 17.185 4.925 ;
      RECT 16.895 4.925 21.025 5.065 ;
      RECT 20.735 5.065 21.025 5.11 ;
      RECT 20.735 4.88 21.025 4.925 ;
      RECT 18.32 1.165 18.64 1.425 ;
      RECT 20.24 1.905 20.56 2.165 ;
      RECT 16.415 4.88 16.705 5.11 ;
      RECT 10.64 5.295 16.63 5.435 ;
      RECT 10.64 5.435 10.96 5.495 ;
      RECT 10.64 5.235 10.96 5.295 ;
      RECT 16.49 5.11 16.63 5.295 ;
      RECT 11.12 5.065 11.44 5.11 ;
      RECT 11.12 4.85 11.44 4.925 ;
      RECT 3.455 4.925 11.44 5.065 ;
      RECT 3.455 5.065 3.745 5.11 ;
      RECT 3.455 4.88 3.745 4.925 ;
      RECT 16.895 1.735 17.185 1.78 ;
      RECT 16.895 1.55 17.185 1.595 ;
      RECT 11.12 1.595 17.185 1.735 ;
      RECT 11.12 1.735 11.44 1.795 ;
      RECT 11.12 1.535 11.44 1.595 ;
      RECT 2.015 5.25 2.305 5.48 ;
      RECT 18.32 5.805 18.64 5.865 ;
      RECT 2.09 5.665 18.64 5.805 ;
      RECT 18.32 5.605 18.64 5.665 ;
      RECT 2.09 5.48 2.23 5.665 ;
      RECT 10.64 1.735 10.96 1.795 ;
      RECT 10.64 1.535 10.96 1.595 ;
      RECT 3.935 1.595 10.96 1.735 ;
      RECT 3.935 1.735 4.225 1.78 ;
      RECT 3.935 1.55 4.225 1.595 ;
  END
END scs8ls_macro_sync_pospos_ret

MACRO scs8ls_macro_sync_sdfrtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.81 2.1 1.265 ;
    END
  END D

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.945 1.44 3.275 2.15 ;
    END
  END SCD

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.26 4.64 1.59 ;
        RECT 3.965 1.18 4.195 1.26 ;
    END
  END CLK

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455 1.66 1.795 1.835 ;
        RECT 0.455 1.49 2.725 1.66 ;
        RECT 2.395 1.26 2.725 1.49 ;
    END
  END SCE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.995 0.35 13.325 1.13 ;
        RECT 13.07 1.13 13.325 2.98 ;
    END
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.44 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.44 3.575 ;
    END
  END vpwr

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3.935 1.965 10.945 2.105 ;
        RECT 3.935 2.105 4.225 2.15 ;
        RECT 7.775 2.105 8.065 2.15 ;
        RECT 10.655 2.105 10.945 2.15 ;
        RECT 3.935 1.92 4.225 1.965 ;
        RECT 7.775 1.92 8.065 1.965 ;
        RECT 10.655 1.92 10.945 1.965 ;
    END
  END RESETB
  OBS
    LAYER mcon ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.995 1.95 4.165 2.12 ;
      RECT 7.835 1.95 8.005 2.12 ;
      RECT 10.715 1.95 10.885 2.12 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
    LAYER li1 ;
      RECT 8.725 1.715 9.005 2.755 ;
      RECT 8.725 1.09 8.895 1.715 ;
      RECT 7.05 0.92 8.895 1.09 ;
      RECT 7.05 1.09 7.325 1.805 ;
      RECT 8.27 0.595 8.655 0.92 ;
      RECT 4.335 1.99 4.585 2.22 ;
      RECT 4.335 1.82 4.98 1.99 ;
      RECT 4.81 1.63 4.98 1.82 ;
      RECT 4.81 1.3 5.28 1.63 ;
      RECT 4.81 1.09 4.98 1.3 ;
      RECT 4.365 0.92 4.98 1.09 ;
      RECT 4.365 0.35 4.535 0.92 ;
      RECT 9.29 2.55 10.315 2.88 ;
      RECT 10.145 1.955 10.315 2.55 ;
      RECT 9.585 1.785 10.315 1.955 ;
      RECT 9.585 1.265 9.755 1.785 ;
      RECT 9.585 1.095 11.395 1.265 ;
      RECT 11.065 1.265 11.395 1.275 ;
      RECT 9.585 0.77 9.755 1.095 ;
      RECT 9.405 0.35 9.755 0.77 ;
      RECT 1.105 0.425 1.435 0.64 ;
      RECT 1.105 0.255 3.605 0.425 ;
      RECT 3.09 0.425 3.605 0.715 ;
      RECT 9.245 2.125 9.975 2.38 ;
      RECT 9.245 1.27 9.415 2.125 ;
      RECT 9.065 0.94 9.415 1.27 ;
      RECT 9.065 0.425 9.235 0.94 ;
      RECT 7.93 0.255 9.235 0.425 ;
      RECT 7.93 0.425 8.1 0.58 ;
      RECT 7.05 0.58 8.1 0.75 ;
      RECT 7.05 0.425 7.22 0.58 ;
      RECT 5.15 0.255 7.22 0.425 ;
      RECT 5.15 0.425 5.62 1.13 ;
      RECT 5.45 1.13 5.62 1.545 ;
      RECT 5.45 1.545 6.2 1.82 ;
      RECT 5.155 1.82 6.2 1.875 ;
      RECT 5.155 1.875 5.62 2.22 ;
      RECT 6.25 2.49 6.88 2.725 ;
      RECT 6.25 2.385 8.075 2.49 ;
      RECT 7.745 2.49 8.075 2.745 ;
      RECT 6.71 2.32 8.075 2.385 ;
      RECT 7.495 1.575 7.665 2.32 ;
      RECT 6.71 1.03 6.88 2.32 ;
      RECT 7.495 1.26 8.315 1.575 ;
      RECT 6.14 0.86 6.88 1.03 ;
      RECT 6.14 0.595 6.47 0.86 ;
      RECT 10.945 2.52 11.31 2.98 ;
      RECT 11.14 1.615 11.31 2.52 ;
      RECT 9.985 1.445 11.735 1.615 ;
      RECT 9.985 1.435 10.315 1.445 ;
      RECT 11.565 0.925 11.735 1.445 ;
      RECT 11.01 0.755 11.735 0.925 ;
      RECT 11.01 0.35 11.34 0.755 ;
      RECT 11.98 2.1 12.31 2.98 ;
      RECT 12.085 1.63 12.31 2.1 ;
      RECT 12.085 1.3 12.87 1.63 ;
      RECT 12.085 0.35 12.335 1.3 ;
      RECT 3.785 1.83 4.165 2.16 ;
      RECT 7.835 1.815 8.165 2.15 ;
      RECT 10.64 1.82 10.97 2.15 ;
      RECT 0.115 2.005 2.705 2.175 ;
      RECT 2.035 1.83 2.705 2.005 ;
      RECT 0.115 2.175 0.445 2.98 ;
      RECT 0.115 1.265 0.285 2.005 ;
      RECT 0.115 0.42 0.365 1.05 ;
      RECT 0.115 1.05 1.375 1.265 ;
      RECT 1.045 0.935 1.375 1.05 ;
      RECT 3.665 2.56 3.995 2.98 ;
      RECT 3.665 2.515 6.075 2.56 ;
      RECT 5.825 2.56 6.075 2.725 ;
      RECT 1.485 2.39 6.075 2.515 ;
      RECT 1.485 2.345 3.995 2.39 ;
      RECT 5.825 2.215 6.075 2.39 ;
      RECT 3.445 2.33 3.995 2.345 ;
      RECT 5.825 2.045 6.54 2.215 ;
      RECT 6.37 1.37 6.54 2.045 ;
      RECT 5.79 1.2 6.54 1.37 ;
      RECT 5.79 0.595 5.96 1.2 ;
      RECT 3.445 1.09 3.615 2.33 ;
      RECT 2.27 0.92 3.615 1.09 ;
      RECT 1.485 2.515 2.555 2.98 ;
      RECT 2.27 0.595 2.6 0.92 ;
      RECT 0 3.245 13.44 3.415 ;
      RECT 4.705 2.73 5.035 3.245 ;
      RECT 3.095 2.685 3.425 3.245 ;
      RECT 7.205 2.66 7.54 3.245 ;
      RECT 10.485 2.52 10.735 3.245 ;
      RECT 11.48 2.1 11.81 3.245 ;
      RECT 12.54 1.82 12.87 3.245 ;
      RECT 8.385 1.745 8.555 3.245 ;
      RECT 0.615 2.345 0.945 3.245 ;
      RECT 0 -0.085 13.44 0.085 ;
      RECT 3.785 0.085 3.955 0.75 ;
      RECT 4.715 0.085 4.965 0.75 ;
      RECT 7.43 0.085 7.76 0.41 ;
      RECT 10.195 0.085 10.525 0.81 ;
      RECT 11.57 0.085 11.905 0.585 ;
      RECT 12.565 0.085 12.815 1.13 ;
      RECT 0.545 0.085 0.875 0.88 ;
  END
END scs8ls_macro_sync_sdfrtp_1

MACRO scs8ls_macro_sync_srsdfrtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 20.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 20.205 0.35 20.535 1.82 ;
        RECT 19.995 1.82 20.535 2.155 ;
        RECT 19.995 2.155 20.325 2.975 ;
    END
  END Q

  PIN RESETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.92 1.55 4.25 1.88 ;
    END
  END RESETB

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.5 0.935 2.17 ;
    END
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.84 2.135 2.17 ;
    END
  END D

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.35 1.55 3.715 1.88 ;
    END
  END SCD

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 16.59 1.46 17.155 1.79 ;
    END
  END CLK

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.235 1.12 18.565 1.45 ;
    END
  END SLEEPB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 20.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 20.64 3.575 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 20.57 2.945 ;
    END
  END kapwr
  OBS
    LAYER mcon ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 15.035 2.735 15.205 2.905 ;
      RECT 15.515 2.735 15.685 2.905 ;
      RECT 17.435 2.735 17.605 2.905 ;
      RECT 15.995 2.735 16.165 2.905 ;
      RECT 20.315 -0.085 20.485 0.085 ;
      RECT 20.315 3.245 20.485 3.415 ;
      RECT 19.835 -0.085 20.005 0.085 ;
      RECT 19.835 3.245 20.005 3.415 ;
      RECT 19.355 -0.085 19.525 0.085 ;
      RECT 19.355 3.245 19.525 3.415 ;
      RECT 18.875 -0.085 19.045 0.085 ;
      RECT 18.875 3.245 19.045 3.415 ;
      RECT 18.395 -0.085 18.565 0.085 ;
      RECT 18.395 3.245 18.565 3.415 ;
      RECT 17.915 -0.085 18.085 0.085 ;
      RECT 17.915 3.245 18.085 3.415 ;
      RECT 17.435 -0.085 17.605 0.085 ;
      RECT 17.435 3.245 17.605 3.415 ;
      RECT 16.955 -0.085 17.125 0.085 ;
      RECT 16.955 2.735 17.125 2.905 ;
      RECT 16.955 3.245 17.125 3.415 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 16.475 2.735 16.645 2.905 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 2.735 14.725 2.905 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
    LAYER li1 ;
      RECT 12.21 2.35 19.325 2.52 ;
      RECT 19.155 1.645 19.325 2.35 ;
      RECT 19.075 1.315 19.345 1.645 ;
      RECT 9.835 2.565 12.54 2.735 ;
      RECT 12.21 2.52 12.54 2.565 ;
      RECT 9.835 2.04 10.5 2.565 ;
      RECT 10.19 0.605 10.5 2.04 ;
      RECT 13.625 2.52 13.955 2.97 ;
      RECT 16.25 1.74 16.42 2.35 ;
      RECT 15.985 1.41 16.42 1.74 ;
      RECT 17.895 1.85 18.49 2.18 ;
      RECT 16.93 0.78 18.345 0.95 ;
      RECT 18.015 0.345 18.345 0.78 ;
      RECT 17.895 0.95 18.065 1.85 ;
      RECT 16.93 0.425 17.1 0.78 ;
      RECT 14.985 0.255 17.1 0.425 ;
      RECT 14.985 0.425 15.315 0.6 ;
      RECT 14.015 0.6 15.315 0.77 ;
      RECT 14.015 0.77 14.185 1.32 ;
      RECT 12.93 1.32 14.185 1.5 ;
      RECT 16.855 2.01 17.495 2.18 ;
      RECT 17.325 1.29 17.495 2.01 ;
      RECT 16.59 1.12 17.495 1.29 ;
      RECT 16.105 1.11 16.76 1.12 ;
      RECT 14.355 0.95 16.76 1.11 ;
      RECT 14.355 1.11 14.525 1.67 ;
      RECT 14.355 0.94 16.435 0.95 ;
      RECT 11.64 1.67 14.525 1.84 ;
      RECT 16.105 0.595 16.435 0.94 ;
      RECT 11.64 1.51 11.97 1.67 ;
      RECT 11.1 2.01 16.08 2.18 ;
      RECT 14.695 1.93 16.08 2.01 ;
      RECT 11.1 1.325 11.43 2.01 ;
      RECT 14.695 1.28 14.955 1.93 ;
      RECT 11.1 1.155 12.235 1.325 ;
      RECT 11.905 0.575 12.235 1.155 ;
      RECT 14.525 2.69 17.73 3.025 ;
      RECT 12.695 0.98 13.845 1.15 ;
      RECT 12.695 0.575 12.945 0.98 ;
      RECT 13.675 0.575 13.845 0.98 ;
      RECT 8.555 2.905 13.455 3.075 ;
      RECT 8.555 2.825 8.725 2.905 ;
      RECT 13.125 2.745 13.455 2.905 ;
      RECT 8.395 2.435 8.725 2.825 ;
      RECT 5.78 2.43 8.725 2.435 ;
      RECT 5.78 2.435 7.68 2.6 ;
      RECT 7.51 2.265 8.725 2.43 ;
      RECT 4.925 2.6 5.95 2.77 ;
      RECT 8.395 1.665 8.725 2.265 ;
      RECT 4.925 1.92 5.095 2.6 ;
      RECT 8.395 1.495 9.4 1.665 ;
      RECT 4.885 1.59 5.215 1.92 ;
      RECT 9.07 1.665 9.4 1.825 ;
      RECT 8.395 1.335 8.99 1.495 ;
      RECT 7.32 1.845 8.135 2.095 ;
      RECT 7.965 1.175 8.135 1.845 ;
      RECT 6.28 1.165 8.135 1.175 ;
      RECT 6.28 1.175 6.61 1.485 ;
      RECT 6.28 1.005 9.53 1.165 ;
      RECT 9.2 1.165 9.53 1.285 ;
      RECT 7.59 0.995 9.53 1.005 ;
      RECT 7.59 0.575 7.84 0.995 ;
      RECT 9.2 0.435 9.53 0.995 ;
      RECT 9.2 0.265 10.93 0.435 ;
      RECT 10.68 0.435 10.93 2.395 ;
      RECT 5.265 2.26 5.555 2.43 ;
      RECT 5.265 2.09 7.11 2.26 ;
      RECT 6.78 1.675 7.11 2.09 ;
      RECT 5.385 1.265 5.555 2.09 ;
      RECT 6.78 1.345 7.795 1.675 ;
      RECT 5.375 0.935 5.555 1.265 ;
      RECT 4.615 0.425 4.865 1.08 ;
      RECT 4.615 0.255 6.59 0.425 ;
      RECT 6.26 0.425 6.59 0.835 ;
      RECT 2.305 2.1 4.755 2.24 ;
      RECT 4.47 2.24 4.755 2.99 ;
      RECT 2.98 2.07 4.715 2.1 ;
      RECT 4.545 1.42 4.715 2.07 ;
      RECT 4.545 1.25 5.205 1.42 ;
      RECT 5.035 0.765 5.205 1.25 ;
      RECT 5.035 0.595 6.055 0.765 ;
      RECT 5.725 0.765 6.055 1.265 ;
      RECT 1.96 2.51 2.635 2.99 ;
      RECT 1.225 2.34 2.635 2.51 ;
      RECT 2.305 2.325 2.635 2.34 ;
      RECT 2.305 2.24 3.08 2.325 ;
      RECT 1.225 1.5 2.08 1.67 ;
      RECT 1.83 0.935 2.08 1.5 ;
      RECT 1.225 1.67 1.395 2.34 ;
      RECT 2.645 1.21 4.375 1.38 ;
      RECT 2.645 0.74 2.975 1.21 ;
      RECT 4.045 0.58 4.375 1.21 ;
      RECT 1.07 0.425 1.32 0.99 ;
      RECT 1.07 0.255 3.405 0.425 ;
      RECT 3.155 0.425 3.405 1.04 ;
      RECT 2.305 1.6 2.88 1.93 ;
      RECT 2.305 0.765 2.475 1.6 ;
      RECT 1.49 0.595 2.475 0.765 ;
      RECT 1.49 0.765 1.66 1.16 ;
      RECT 0.105 1.16 1.66 1.33 ;
      RECT 0.105 1.33 0.435 2.99 ;
      RECT 0.105 0.53 0.355 1.16 ;
      RECT 0 -0.085 20.64 0.085 ;
      RECT 18.805 0.085 19.055 0.805 ;
      RECT 19.855 0.085 20.025 1.13 ;
      RECT 0.535 0.085 0.865 0.99 ;
      RECT 3.615 0.085 3.865 1.04 ;
      RECT 7.05 0.085 7.38 0.835 ;
      RECT 8.02 0.085 8.35 0.825 ;
      RECT 11.365 0.085 11.695 0.985 ;
      RECT 13.125 0.085 13.455 0.81 ;
      RECT 17.475 0.085 17.805 0.61 ;
      RECT 0 3.245 20.64 3.415 ;
      RECT 6.12 2.77 6.45 3.245 ;
      RECT 7.85 2.605 8.18 3.245 ;
      RECT 3.245 2.41 4.3 3.245 ;
      RECT 19.495 1.815 19.825 3.245 ;
      RECT 0.645 2.34 0.975 3.245 ;
      RECT 19.515 1.315 20.02 1.645 ;
      RECT 18.735 1.815 18.985 2.18 ;
      RECT 18.735 1.145 18.905 1.815 ;
      RECT 18.735 0.975 19.685 1.145 ;
      RECT 19.515 1.145 19.685 1.315 ;
      RECT 19.235 0.345 19.685 0.975 ;
  END
END scs8ls_macro_sync_srsdfrtp_1

MACRO scs8ls_macro_sparecell
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 13.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.92 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.92 0.245 ;
    END
  END vgnd

  PIN LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.415 1.58 9.505 1.75 ;
        RECT 4.415 1.75 4.705 1.78 ;
        RECT 5.375 1.75 5.665 1.78 ;
        RECT 7.295 1.75 7.585 1.78 ;
        RECT 8.255 1.75 8.545 1.78 ;
        RECT 9.215 1.75 9.505 1.78 ;
        RECT 4.415 1.55 4.705 1.58 ;
        RECT 5.375 1.55 5.665 1.58 ;
        RECT 7.295 1.55 7.585 1.58 ;
        RECT 8.255 1.55 8.545 1.58 ;
        RECT 9.215 1.55 9.505 1.58 ;
    END
    ANTENNADIFFAREA 2.3828 ;
    ANTENNAGATEAREA 2.232 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 3.654 LAYER met1 ;
  END LO

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 13.115 1.21 13.285 1.38 ;
      RECT 13.115 1.58 13.285 1.75 ;
      RECT 12.635 1.58 12.805 1.75 ;
      RECT 12.155 1.21 12.325 1.38 ;
      RECT 10.715 1.58 10.885 1.75 ;
      RECT 10.235 1.21 10.405 1.38 ;
      RECT 9.755 1.21 9.925 1.38 ;
      RECT 9.275 1.58 9.445 1.75 ;
      RECT 8.315 1.58 8.485 1.75 ;
      RECT 7.355 1.58 7.525 1.75 ;
      RECT 5.435 1.58 5.605 1.75 ;
      RECT 4.475 1.58 4.645 1.75 ;
      RECT 3.995 1.21 4.165 1.38 ;
      RECT 3.515 1.21 3.685 1.38 ;
      RECT 3.035 1.58 3.205 1.75 ;
      RECT 1.595 1.21 1.765 1.38 ;
      RECT 1.115 1.58 1.285 1.75 ;
      RECT 0.635 1.21 0.805 1.38 ;
      RECT 0.635 1.58 0.805 1.75 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
    LAYER met1 ;
      RECT 13.055 1.18 13.345 1.78 ;
      RECT 10.655 1.75 10.945 1.78 ;
      RECT 10.655 1.58 12.865 1.75 ;
      RECT 12.575 1.75 12.865 1.78 ;
      RECT 10.655 1.55 10.945 1.58 ;
      RECT 12.575 1.55 12.865 1.58 ;
      RECT 9.695 1.38 9.985 1.41 ;
      RECT 9.695 1.21 12.385 1.38 ;
      RECT 10.175 1.38 10.465 1.41 ;
      RECT 12.095 1.38 12.385 1.41 ;
      RECT 9.695 1.18 9.985 1.21 ;
      RECT 10.175 1.18 10.465 1.21 ;
      RECT 12.095 1.18 12.385 1.21 ;
      RECT 1.535 1.38 1.825 1.41 ;
      RECT 1.535 1.21 4.225 1.38 ;
      RECT 3.455 1.38 3.745 1.41 ;
      RECT 3.935 1.38 4.225 1.41 ;
      RECT 1.535 1.18 1.825 1.21 ;
      RECT 3.455 1.18 3.745 1.21 ;
      RECT 3.935 1.18 4.225 1.21 ;
      RECT 1.055 1.75 1.345 1.78 ;
      RECT 1.055 1.58 3.265 1.75 ;
      RECT 2.975 1.75 3.265 1.78 ;
      RECT 1.055 1.55 1.345 1.58 ;
      RECT 2.975 1.55 3.265 1.58 ;
      RECT 0.575 1.18 0.865 1.78 ;
    LAYER li1 ;
      RECT 1.565 0.44 2.035 1.41 ;
      RECT 1.705 1.41 2.035 1.605 ;
      RECT 1.705 0.255 2.035 0.44 ;
      RECT 11.885 0.44 12.355 1.41 ;
      RECT 11.885 1.41 12.215 1.605 ;
      RECT 11.885 0.255 12.215 0.44 ;
      RECT 2.895 1.82 3.235 2.735 ;
      RECT 2.895 0.35 3.225 1.82 ;
      RECT 10.685 1.82 11.025 2.735 ;
      RECT 10.695 0.35 11.025 1.82 ;
      RECT 3.395 1.18 3.725 1.55 ;
      RECT 10.195 1.18 10.525 1.55 ;
      RECT 1.555 1.945 1.885 2.98 ;
      RECT 1.555 1.775 2.705 1.945 ;
      RECT 2.535 1.945 2.705 2.905 ;
      RECT 2.535 2.905 3.685 3.075 ;
      RECT 3.435 1.82 3.685 2.905 ;
      RECT 10.235 2.905 11.385 3.075 ;
      RECT 11.215 1.945 11.385 2.905 ;
      RECT 10.235 1.82 10.485 2.905 ;
      RECT 11.215 1.775 12.365 1.945 ;
      RECT 12.035 1.945 12.365 2.98 ;
      RECT 2.085 2.115 2.335 3.245 ;
      RECT 3.98 2.29 4.31 3.245 ;
      RECT 4.89 2.29 5.22 3.245 ;
      RECT 5.87 1.82 6.12 3.245 ;
      RECT 1.005 1.95 1.335 3.245 ;
      RECT 0.105 1.82 0.355 3.245 ;
      RECT 6.525 2.505 6.855 3.245 ;
      RECT 8.7 2.29 9.03 3.245 ;
      RECT 9.61 2.29 9.94 3.245 ;
      RECT 7.8 1.82 8.05 3.245 ;
      RECT 11.585 2.115 11.835 3.245 ;
      RECT 12.585 1.95 12.915 3.245 ;
      RECT 13.565 1.82 13.815 3.245 ;
      RECT 0 3.245 13.92 3.415 ;
      RECT 2.395 0.085 2.725 1.13 ;
      RECT 3.395 0.085 3.725 1.01 ;
      RECT 5.365 0.085 5.695 0.84 ;
      RECT 0.12 0.085 0.37 1.13 ;
      RECT 1.06 0.085 1.31 1.13 ;
      RECT 7.065 0.085 7.395 0.825 ;
      RECT 8.225 0.085 8.555 0.84 ;
      RECT 10.195 0.085 10.525 1.01 ;
      RECT 11.195 0.085 11.525 1.13 ;
      RECT 12.61 0.085 12.86 1.13 ;
      RECT 13.55 0.085 13.8 1.13 ;
      RECT 0 -0.085 13.92 0.085 ;
      RECT 4.425 1.35 4.755 1.78 ;
      RECT 9.165 1.35 9.495 1.78 ;
      RECT 4.925 1.35 5.635 1.78 ;
      RECT 8.285 1.35 8.995 1.78 ;
      RECT 3.965 1.18 4.195 1.95 ;
      RECT 3.965 1.95 5.67 2.12 ;
      RECT 3.965 1.01 4.785 1.18 ;
      RECT 4.51 2.12 4.68 2.98 ;
      RECT 5.42 2.12 5.67 2.98 ;
      RECT 4.455 0.595 4.785 1.01 ;
      RECT 9.725 1.18 9.955 1.95 ;
      RECT 8.25 1.95 9.955 2.12 ;
      RECT 9.135 1.01 9.955 1.18 ;
      RECT 8.25 2.12 8.5 2.98 ;
      RECT 9.24 2.12 9.41 2.98 ;
      RECT 9.135 0.595 9.465 1.01 ;
      RECT 4.965 1.01 6.125 1.18 ;
      RECT 4.965 0.425 5.135 1.01 ;
      RECT 5.875 0.35 6.125 1.01 ;
      RECT 3.955 0.255 5.135 0.425 ;
      RECT 3.955 0.425 4.285 0.84 ;
      RECT 7.795 1.01 8.955 1.18 ;
      RECT 8.785 0.425 8.955 1.01 ;
      RECT 7.795 0.35 8.045 1.01 ;
      RECT 8.785 0.255 9.965 0.425 ;
      RECT 9.635 0.425 9.965 0.84 ;
      RECT 13.085 1.13 13.37 2.98 ;
      RECT 13.04 0.35 13.37 1.13 ;
      RECT 0.55 1.13 0.835 2.98 ;
      RECT 0.55 0.35 0.88 1.13 ;
      RECT 1.005 1.3 1.335 1.78 ;
      RECT 12.585 1.3 12.915 1.78 ;
      RECT 7.295 0.995 7.595 2.485 ;
      RECT 7.065 2.485 7.595 3.075 ;
      RECT 6.325 0.845 6.635 2.335 ;
      RECT 6.325 0.255 6.855 0.845 ;
  END
END scs8ls_macro_sparecell
  
END LIBRARY
