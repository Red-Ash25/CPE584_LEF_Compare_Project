# 
# LEF OUT 
# User Name : iptguser 
# Date : Mon Feb  4 15:39:14 2013
# 
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO scs8ls_lpflow_decaphekapwr_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.96 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 0.89 2.945 ;
    END
  END kapwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.96 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 0.96 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 0.96 3.415 ;
      RECT 0.085 0.085 0.47 1.675 ;
      RECT 0 -0.085 0.96 0.085 ;
      RECT 0.085 1.845 0.875 3.075 ;
    LAYER mcon ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.575 2.725 0.745 2.895 ;
      RECT 0.215 2.725 0.385 2.895 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_lpflow_decaphekapwr_2

MACRO scs8ls_lpflow_decaphekapwr_3
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
    END
  END vgnd

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 1.37 2.945 ;
    END
  END kapwr

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 1.44 3.415 ;
      RECT 0.085 1.77 1.355 3.075 ;
      RECT 0.805 1.25 1.355 1.77 ;
      RECT 0.085 1.08 0.635 1.6 ;
      RECT 0.085 0.085 1.355 1.08 ;
      RECT 0 -0.085 1.44 0.085 ;
    LAYER mcon ;
      RECT 0.85 2.725 1.02 2.895 ;
      RECT 0.42 2.725 0.59 2.895 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_decaphekapwr_3

MACRO scs8ls_lpflow_decaphekapwr_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 1.85 2.945 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 1.92 3.415 ;
      RECT 0.085 1.77 1.835 3.075 ;
      RECT 1.06 1.25 1.835 1.77 ;
      RECT 0.085 1.08 0.89 1.6 ;
      RECT 0.085 0.085 1.835 1.08 ;
      RECT 0 -0.085 1.92 0.085 ;
    LAYER mcon ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.49 2.725 0.66 2.895 ;
      RECT 0.85 2.725 1.02 2.895 ;
      RECT 1.21 2.725 1.38 2.895 ;
  END
END scs8ls_lpflow_decaphekapwr_4

MACRO scs8ls_lpflow_decaphekapwr_6
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 2.81 2.945 ;
    END
  END kapwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.085 1.77 2.795 3.075 ;
      RECT 1.365 1.25 2.795 1.77 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 0.085 1.08 1.195 1.6 ;
      RECT 0.085 0.085 2.795 1.08 ;
      RECT 0 -0.085 2.88 0.085 ;
    LAYER mcon ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.895 2.725 2.065 2.895 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 0.815 2.725 0.985 2.895 ;
      RECT 2.255 2.725 2.425 2.895 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 0.455 2.725 0.625 2.895 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 1.535 2.725 1.705 2.895 ;
      RECT 1.175 2.725 1.345 2.895 ;
  END
END scs8ls_lpflow_decaphekapwr_6

MACRO scs8ls_lpflow_decaphekapwr_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 3.77 2.945 ;
    END
  END kapwr

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.085 1.075 0.95 1.6 ;
      RECT 0.085 1.07 2.71 1.075 ;
      RECT 2 1.075 2.71 1.6 ;
      RECT 0.085 0.085 3.755 1.07 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 0.085 1.77 3.755 3.075 ;
      RECT 1.12 1.25 1.83 1.77 ;
      RECT 2.88 1.25 3.755 1.77 ;
      RECT 0 3.245 3.84 3.415 ;
    LAYER mcon ;
      RECT 0.49 2.725 0.66 2.895 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 1.21 2.725 1.38 2.895 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 2.34 2.725 2.51 2.895 ;
      RECT 3.06 2.725 3.23 2.895 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.7 2.725 2.87 2.895 ;
      RECT 1.62 2.725 1.79 2.895 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 1.98 2.725 2.15 2.895 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.85 2.725 1.02 2.895 ;
      RECT 2.075 3.245 2.245 3.415 ;
  END
END scs8ls_lpflow_decaphekapwr_8

MACRO scs8ls_lpflow_inputiso0n_lp
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY R90 ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.345 1.395 1.09 1.75 ;
    END
    ANTENNAGATEAREA 0.189 LAYER met1 ;
    ANTENNAGATEAREA 0.189 LAYER met2 ;
    ANTENNAGATEAREA 0.189 LAYER met3 ;
    ANTENNAGATEAREA 0.189 LAYER met4 ;
    ANTENNAGATEAREA 0.189 LAYER met5 ;
  END A

  PIN sleepb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.315 1.395 1.985 1.75 ;
    END
    ANTENNAGATEAREA 0.189 LAYER met1 ;
    ANTENNAGATEAREA 0.189 LAYER met2 ;
    ANTENNAGATEAREA 0.189 LAYER met3 ;
    ANTENNAGATEAREA 0.189 LAYER met4 ;
    ANTENNAGATEAREA 0.189 LAYER met5 ;
  END sleepb

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855 0.465 3.275 3.075 ;
    END
    ANTENNADIFFAREA 0.4081 LAYER met1 ;
    ANTENNADIFFAREA 0.4081 LAYER met2 ;
    ANTENNADIFFAREA 0.4081 LAYER met3 ;
    ANTENNADIFFAREA 0.4081 LAYER met4 ;
    ANTENNADIFFAREA 0.4081 LAYER met5 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 1.44 0.085 2.335 0.84 ;
      RECT 1.08 2.125 1.41 2.82 ;
      RECT 1.08 1.955 2.685 2.125 ;
      RECT 2.275 1.225 2.685 1.955 ;
      RECT 0.65 1.055 2.685 1.225 ;
      RECT 0.65 0.51 0.98 1.055 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 0.29 2.345 0.62 3.245 ;
      RECT 1.99 2.295 2.675 3.245 ;
    LAYER mcon ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_inputiso0n_lp

MACRO scs8ls_lpflow_inputiso0n_lp2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY R90 ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045 0.765 2.275 2.015 ;
        RECT 1.795 2.015 2.275 3.065 ;
        RECT 1.945 0.305 2.275 0.765 ;
    END
    ANTENNADIFFAREA 0.4047 LAYER met1 ;
    ANTENNADIFFAREA 0.4047 LAYER met2 ;
    ANTENNADIFFAREA 0.4047 LAYER met3 ;
    ANTENNADIFFAREA 0.4047 LAYER met4 ;
    ANTENNADIFFAREA 0.4047 LAYER met5 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.955 0.455 1.78 ;
    END
    ANTENNAGATEAREA 0.313 LAYER met1 ;
    ANTENNAGATEAREA 0.313 LAYER met2 ;
    ANTENNAGATEAREA 0.313 LAYER met3 ;
    ANTENNAGATEAREA 0.313 LAYER met4 ;
    ANTENNAGATEAREA 0.313 LAYER met5 ;
  END A

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1 1.515 1.795 1.845 ;
        RECT 1 1.445 1.33 1.515 ;
    END
    ANTENNAGATEAREA 0.313 LAYER met1 ;
    ANTENNAGATEAREA 0.313 LAYER met2 ;
    ANTENNAGATEAREA 0.313 LAYER met3 ;
    ANTENNAGATEAREA 0.313 LAYER met4 ;
    ANTENNAGATEAREA 0.313 LAYER met5 ;
  END SLEEPB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.65 0.945 1.81 1.275 ;
      RECT 0.65 2.015 1.065 3.065 ;
      RECT 0.65 1.275 0.82 2.015 ;
      RECT 0.65 0.765 0.82 0.945 ;
      RECT 0.305 0.595 0.82 0.765 ;
      RECT 0.305 0.305 0.635 0.595 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 1.085 0.085 1.455 0.765 ;
      RECT 0 3.245 2.4 3.415 ;
      RECT 0.14 2.015 0.47 3.245 ;
      RECT 1.265 2.015 1.595 3.245 ;
    LAYER mcon ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
  END
END scs8ls_lpflow_inputiso0n_lp2

MACRO scs8ls_lpflow_inputiso0p_lp
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY R90 ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.98 1.395 2.65 1.75 ;
    END
    ANTENNAGATEAREA 0.189 LAYER met1 ;
    ANTENNAGATEAREA 0.189 LAYER met2 ;
    ANTENNAGATEAREA 0.189 LAYER met3 ;
    ANTENNAGATEAREA 0.189 LAYER met4 ;
    ANTENNAGATEAREA 0.189 LAYER met5 ;
  END A

  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.16 0.92 1.895 ;
    END
    ANTENNAGATEAREA 0.252 LAYER met1 ;
    ANTENNAGATEAREA 0.252 LAYER met2 ;
    ANTENNAGATEAREA 0.252 LAYER met3 ;
    ANTENNAGATEAREA 0.252 LAYER met4 ;
    ANTENNAGATEAREA 0.252 LAYER met5 ;
  END sleep

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.4 0.465 3.755 3.075 ;
    END
    ANTENNADIFFAREA 0.4081 LAYER met1 ;
    ANTENNADIFFAREA 0.4081 LAYER met2 ;
    ANTENNADIFFAREA 0.4081 LAYER met3 ;
    ANTENNADIFFAREA 0.4081 LAYER met4 ;
    ANTENNADIFFAREA 0.4081 LAYER met5 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.155 2.065 1.595 2.235 ;
      RECT 1.2 1.39 1.595 2.065 ;
      RECT 0.155 2.235 0.375 2.855 ;
      RECT 0.155 0.43 0.375 2.065 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 0.895 2.41 1.225 3.245 ;
      RECT 2.525 2.295 2.91 3.245 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 0.895 0.085 1.575 0.84 ;
      RECT 2.55 0.085 2.885 0.835 ;
      RECT 1.765 1.955 3.23 2.125 ;
      RECT 2.82 1.225 3.23 1.955 ;
      RECT 2.095 1.005 3.23 1.225 ;
      RECT 2.095 0.43 2.305 1.005 ;
      RECT 1.765 2.125 1.975 2.855 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_inputiso0p_lp

MACRO scs8ls_lpflow_inputiso0p_lp2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY R90 ;
  SITE unit ;

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.01 0.92 1.78 ;
    END
    ANTENNAGATEAREA 0.376 LAYER met1 ;
    ANTENNAGATEAREA 0.376 LAYER met2 ;
    ANTENNAGATEAREA 0.376 LAYER met3 ;
    ANTENNAGATEAREA 0.376 LAYER met4 ;
    ANTENNAGATEAREA 0.376 LAYER met5 ;
  END SLEEP

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.4 0.465 3.755 3.075 ;
    END
    ANTENNADIFFAREA 0.3763 LAYER met1 ;
    ANTENNADIFFAREA 0.3763 LAYER met2 ;
    ANTENNADIFFAREA 0.3763 LAYER met3 ;
    ANTENNADIFFAREA 0.3763 LAYER met4 ;
    ANTENNADIFFAREA 0.3763 LAYER met5 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.98 1.395 2.755 1.75 ;
    END
    ANTENNAGATEAREA 0.313 LAYER met1 ;
    ANTENNAGATEAREA 0.313 LAYER met2 ;
    ANTENNAGATEAREA 0.313 LAYER met3 ;
    ANTENNAGATEAREA 0.313 LAYER met4 ;
    ANTENNAGATEAREA 0.313 LAYER met5 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 2.235 2.295 3.145 3.245 ;
      RECT 0.635 2.29 1.485 3.245 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 0.895 0.085 1.575 0.84 ;
      RECT 2.55 0.085 2.885 0.835 ;
      RECT 1.765 1.955 3.23 2.125 ;
      RECT 2.925 1.225 3.23 1.955 ;
      RECT 2.095 1.005 3.23 1.225 ;
      RECT 2.095 0.43 2.305 1.005 ;
      RECT 1.765 2.125 1.975 3.075 ;
      RECT 0.155 1.95 1.595 2.12 ;
      RECT 1.2 1.01 1.595 1.95 ;
      RECT 0.155 2.12 0.375 3.075 ;
      RECT 0.155 0.43 0.375 1.95 ;
    LAYER mcon ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_inputiso0p_lp2

MACRO scs8ls_lpflow_inputiso1n_lp
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.91 1.395 2.58 1.75 ;
    END
    ANTENNAGATEAREA 0.189 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.137 LAYER li1 ;
  END A

  PIN sleepb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.54 1.16 1.16 1.99 ;
    END
    ANTENNAGATEAREA 0.252 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.154 LAYER li1 ;
  END sleepb

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395 0.465 3.755 3.075 ;
    END
    ANTENNADIFFAREA 0.4081 ;
    ANTENNAPARTIALMETALSIDEAREA 0.254 LAYER li1 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.095 2.125 2.305 2.88 ;
      RECT 2.095 1.955 3.225 2.125 ;
      RECT 2.895 1.225 3.225 1.955 ;
      RECT 1.87 1.055 3.225 1.225 ;
      RECT 1.87 0.885 2.065 1.055 ;
      RECT 1.735 0.43 2.065 0.885 ;
      RECT 0.345 2.33 0.59 2.82 ;
      RECT 0.125 2.16 1.7 2.33 ;
      RECT 1.37 1.315 1.7 2.16 ;
      RECT 0.125 0.885 0.37 2.16 ;
      RECT 0.12 0.43 0.365 0.885 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 0.885 0.085 1.215 0.885 ;
      RECT 2.525 0.085 2.855 0.885 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 1.19 2.5 1.52 3.245 ;
      RECT 2.525 2.295 2.91 3.245 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_inputiso1n_lp

MACRO scs8ls_lpflow_inputiso1p_lp
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435 1.35 2.105 1.75 ;
    END
    ANTENNAGATEAREA 0.189 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.146 LAYER li1 ;
  END sleep

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855 0.465 3.275 3.075 ;
    END
    ANTENNADIFFAREA 0.4081 ;
    ANTENNAPARTIALMETALSIDEAREA 0.266 LAYER li1 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555 1.16 0.855 1.35 ;
        RECT 0.555 1.35 1.225 1.75 ;
    END
    ANTENNAGATEAREA 0.189 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.116 LAYER li1 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 1.56 2.295 2.365 3.245 ;
      RECT 0.77 1.955 2.685 2.125 ;
      RECT 2.35 1.18 2.685 1.955 ;
      RECT 1.28 1.01 2.685 1.18 ;
      RECT 1.28 0.44 1.49 1.01 ;
      RECT 0.77 2.125 1.1 2.82 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 0.46 0.085 0.76 0.84 ;
      RECT 2.01 0.085 2.34 0.84 ;
    LAYER mcon ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_inputiso1p_lp

MACRO scs8ls_lpflow_inputisolatch_lp
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SLEEPB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.585 1.455 5.255 1.785 ;
    END
    ANTENNAGATEAREA 0.222 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.132 LAYER li1 ;
  END SLEEPB

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.755 0.44 7.085 2.955 ;
    END
    ANTENNADIFFAREA 0.4047 ;
    ANTENNAPARTIALMETALSIDEAREA 0.229 LAYER li1 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.465 1.185 1.27 1.78 ;
        RECT 0.465 1.78 0.825 2.755 ;
    END
    ANTENNAGATEAREA 0.126 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.339 LAYER li1 ;
  END D

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 5.445 0.43 5.875 0.745 ;
      RECT 4.045 1.955 6.025 2.125 ;
      RECT 5.695 2.125 6.025 2.955 ;
      RECT 5.695 1.915 6.025 1.955 ;
      RECT 5.705 0.745 5.875 1.915 ;
      RECT 4.045 1.505 4.375 1.955 ;
      RECT 3.705 2.295 4.985 2.465 ;
      RECT 4.045 2.465 4.985 2.975 ;
      RECT 2.24 1.335 2.49 1.455 ;
      RECT 2.24 1.165 4.035 1.335 ;
      RECT 2.24 1.125 2.49 1.165 ;
      RECT 3.865 0.845 4.035 1.165 ;
      RECT 3.705 1.335 3.875 2.295 ;
      RECT 3.865 0.595 4.195 0.845 ;
      RECT 1.445 2.805 2.41 2.975 ;
      RECT 1.445 1.795 1.615 2.805 ;
      RECT 2.24 1.795 2.41 2.805 ;
      RECT 1.445 1.125 1.73 1.795 ;
      RECT 2.24 1.625 3.535 1.795 ;
      RECT 1.445 1.015 1.615 1.125 ;
      RECT 3.285 1.795 3.535 3 ;
      RECT 0.16 0.845 1.615 1.015 ;
      RECT 0.16 0.375 0.41 0.845 ;
      RECT 4.365 0.845 5.115 0.915 ;
      RECT 4.365 0.915 5.535 1.015 ;
      RECT 4.945 1.015 5.535 1.245 ;
      RECT 1.795 1.965 2.07 2.635 ;
      RECT 1.9 0.955 2.07 1.965 ;
      RECT 1.785 0.825 3.695 0.955 ;
      RECT 2.63 0.955 3.695 0.995 ;
      RECT 1.785 0.785 2.8 0.825 ;
      RECT 3.525 0.425 3.695 0.825 ;
      RECT 1.785 0.325 2.285 0.785 ;
      RECT 3.525 0.255 4.535 0.425 ;
      RECT 4.365 0.425 4.535 0.845 ;
      RECT 0 -0.085 7.2 0.085 ;
      RECT 0.59 0.085 0.92 0.675 ;
      RECT 3.105 0.085 3.355 0.655 ;
      RECT 4.705 0.085 4.985 0.675 ;
      RECT 6.045 0.085 6.295 1.26 ;
      RECT 0 3.245 7.2 3.415 ;
      RECT 0.995 2.54 1.265 3.245 ;
      RECT 5.155 2.295 5.485 3.245 ;
      RECT 2.755 1.965 3.085 3.245 ;
      RECT 6.225 1.915 6.555 3.245 ;
    LAYER mcon ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
  END
END scs8ls_lpflow_inputisolatch_lp

MACRO scs8ls_lpflow_lsbuf_hl_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.515 0.35 2.765 1.35 ;
        RECT 1.755 1.35 2.765 1.6 ;
        RECT 2.515 1.6 2.765 2.98 ;
        RECT 1.755 1.6 1.925 1.82 ;
        RECT 1.755 1.13 1.925 1.35 ;
        RECT 1.595 1.82 1.925 2.98 ;
        RECT 1.685 0.35 1.925 1.13 ;
    END
    ANTENNADIFFAREA 1.0864 ;
    ANTENNAPARTIALMETALSIDEAREA 1.114 LAYER li1 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.45 0.905 1.78 ;
    END
    ANTENNAGATEAREA 0.363 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.09 LAYER li1 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN lowlvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 3.29 2.945 ;
    END
  END lowlvpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.935 0.085 3.205 1.13 ;
      RECT 0.76 0.085 1.515 0.94 ;
      RECT 2.095 0.085 2.345 1.13 ;
      RECT 0.12 2.1 0.4 2.98 ;
      RECT 2.935 1.82 3.255 2.98 ;
      RECT 2.095 1.82 2.345 2.98 ;
      RECT 1.095 2.29 1.425 2.98 ;
      RECT 0.57 2.12 0.875 2.98 ;
      RECT 0.57 1.95 1.245 2.12 ;
      RECT 1.075 1.63 1.245 1.95 ;
      RECT 1.075 1.3 1.585 1.63 ;
      RECT 1.075 1.28 1.245 1.3 ;
      RECT 0.33 1.11 1.245 1.28 ;
      RECT 0.33 0.35 0.59 1.11 ;
      RECT 0 3.245 3.36 3.415 ;
    LAYER mcon ;
      RECT 0.175 2.73 0.345 2.9 ;
      RECT 3.005 2.73 3.175 2.9 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.135 2.73 2.305 2.9 ;
      RECT 1.175 2.73 1.345 2.9 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
  END
END scs8ls_lpflow_lsbuf_hl_4

MACRO scs8ls_lpflow_lsbuf_hl_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.47 1.82 1.8 2.98 ;
        RECT 1.63 1.13 1.8 1.82 ;
        RECT 1.475 0.35 1.8 1.13 ;
    END
    ANTENNADIFFAREA 0.5432 ;
    ANTENNAPARTIALMETALSIDEAREA 0.419 LAYER li1 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.45 0.91 1.78 ;
    END
    ANTENNAGATEAREA 0.2085 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.087 LAYER li1 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN lowlvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 2.33 2.945 ;
    END
  END lowlvpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.97 1.82 2.25 2.98 ;
      RECT 0.97 2.29 1.3 2.98 ;
      RECT 0.47 2.12 0.8 2.98 ;
      RECT 0.47 1.95 1.3 2.12 ;
      RECT 1.13 1.63 1.3 1.95 ;
      RECT 1.13 1.3 1.46 1.63 ;
      RECT 1.13 1.28 1.3 1.3 ;
      RECT 0.115 1.11 1.3 1.28 ;
      RECT 0.115 0.8 0.795 1.11 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 1.97 0.085 2.235 1.13 ;
      RECT 0.975 0.085 1.305 0.94 ;
      RECT 0 3.245 2.4 3.415 ;
    LAYER mcon ;
      RECT 2 2.73 2.17 2.9 ;
      RECT 1.05 2.73 1.22 2.9 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
  END
END scs8ls_lpflow_lsbuf_hl_2

MACRO scs8ls_lpflow_lsbuf_hl_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.47 1.82 1.83 2.98 ;
        RECT 1.66 1.13 1.83 1.82 ;
        RECT 1.475 0.35 1.83 1.13 ;
    END
    ANTENNADIFFAREA 0.5413 ;
    ANTENNAPARTIALMETALSIDEAREA 0.431 LAYER li1 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.45 0.91 1.78 ;
    END
    ANTENNAGATEAREA 0.2085 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.087 LAYER li1 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr

  PIN lowlvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 1.85 2.945 ;
    END
  END lowlvpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.97 2.29 1.3 2.98 ;
      RECT 1.13 1.3 1.49 1.63 ;
      RECT 0.47 2.12 0.8 2.98 ;
      RECT 0.47 1.95 1.3 2.12 ;
      RECT 1.13 1.63 1.3 1.95 ;
      RECT 1.13 1.28 1.3 1.3 ;
      RECT 0.115 1.11 1.3 1.28 ;
      RECT 0.115 0.8 0.795 1.11 ;
      RECT 0 -0.085 1.92 0.085 ;
      RECT 0.975 0.085 1.305 0.94 ;
      RECT 0 3.245 1.92 3.415 ;
    LAYER mcon ;
      RECT 1.05 2.73 1.22 2.9 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_lsbuf_hl_1

MACRO scs8ls_lpflow_lsbuf_lh_isowell_tap_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.59 6.595 2.98 ;
        RECT 5.465 1.36 6.595 1.59 ;
        RECT 5.465 1.59 5.695 2.98 ;
        RECT 5.465 0.35 5.695 1.36 ;
        RECT 6.365 0.35 6.595 1.36 ;
    END
    ANTENNADIFFAREA 1.0864 ;
    ANTENNAPARTIALMETALSIDEAREA 1.096 LAYER li1 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.83 3.29 2.15 ;
        RECT 2.97 1.56 3.63 1.83 ;
        RECT 2.97 1.5 3.445 1.56 ;
    END
    ANTENNAGATEAREA 0.675 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER li1 ;
  END A

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 4.125 7.13 4.385 ;
    END
  END vpb

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
    END
  END vpwr

  PIN lowlvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 7.13 2.945 ;
    END
  END lowlvpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 7.2 6.905 ;
    END
  END vgnd
  OBS
    LAYER li1 ;
      RECT 6.895 5.59 7.065 6.575 ;
      RECT 0 6.575 7.2 6.745 ;
      RECT 4.365 5.53 5.035 6.575 ;
      RECT 3.505 5.53 3.835 6.575 ;
      RECT 2.645 5.53 2.975 6.575 ;
      RECT 0.135 5.59 0.305 6.575 ;
      RECT 0 -0.085 7.2 0.085 ;
      RECT 6.765 0.085 7.075 1.13 ;
      RECT 0.135 0.085 0.305 1.07 ;
      RECT 3.115 0.085 3.445 1.13 ;
      RECT 3.975 0.085 4.305 1.05 ;
      RECT 4.91 0.085 5.24 1.13 ;
      RECT 2.02 0.085 2.35 1.13 ;
      RECT 5.865 0.085 6.195 1.13 ;
      RECT 6.87 3.65 7.1 4.4 ;
      RECT 0.1 3.65 0.33 4.4 ;
      RECT 6.765 1.82 7.095 3.245 ;
      RECT 4.89 3.245 7.2 3.415 ;
      RECT 4.89 1.82 5.235 3.245 ;
      RECT 4.89 3.415 5.12 4.84 ;
      RECT 5.865 1.82 6.195 3.245 ;
      RECT 3.615 1.22 4.665 1.39 ;
      RECT 3.615 0.35 3.805 1.22 ;
      RECT 4.475 0.35 4.665 1.22 ;
      RECT 3.68 3.185 3.85 4.235 ;
      RECT 3.68 3.015 4.19 3.185 ;
      RECT 4.02 1.39 4.19 3.015 ;
      RECT 4.39 4.405 4.72 4.84 ;
      RECT 3.68 4.235 4.72 4.405 ;
      RECT 4.39 3.695 4.72 4.235 ;
      RECT 3.145 5.19 5.19 5.36 ;
      RECT 4.6 5.01 5.19 5.19 ;
      RECT 4.005 5.36 4.195 6.31 ;
      RECT 3.145 5.36 3.335 6.31 ;
      RECT 5.205 5.53 5.55 6.31 ;
      RECT 5.36 3.915 5.55 5.53 ;
      RECT 5.36 3.585 6.41 3.915 ;
      RECT 3.06 4.77 3.73 5.02 ;
      RECT 3.06 2.98 3.3 4.77 ;
      RECT 2.56 2.74 3.3 2.98 ;
      RECT 2.56 0.735 2.8 2.74 ;
      RECT 0 3.245 1.89 3.415 ;
      RECT 4.02 3.525 4.19 4.065 ;
      RECT 4.02 3.355 4.64 3.525 ;
      RECT 4.47 1.82 4.64 3.355 ;
      RECT 2.06 3.27 2.81 3.94 ;
      RECT 2.06 2.945 2.39 3.27 ;
      RECT 1.38 2.675 2.39 2.945 ;
      RECT 2.06 1.9 2.39 2.675 ;
    LAYER mcon ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.14 2.715 2.31 2.885 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 6.9 4.17 7.07 4.34 ;
      RECT 0.13 4.17 0.3 4.34 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 6.395 6.575 6.565 6.745 ;
      RECT 6.875 6.575 7.045 6.745 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 1.42 2.725 1.59 2.895 ;
      RECT 1.78 2.725 1.95 2.895 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 3.035 6.575 3.205 6.745 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
  END
END scs8ls_lpflow_lsbuf_lh_isowell_tap_4

MACRO scs8ls_lpflow_lsbuf_lh_isowell_tap_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.24 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.355 1.3 5.685 2.98 ;
        RECT 5.355 0.35 5.59 1.3 ;
    END
    ANTENNADIFFAREA 0.5432 ;
    ANTENNAPARTIALMETALSIDEAREA 0.456 LAYER li1 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.83 3.29 2.15 ;
        RECT 2.97 1.56 3.63 1.83 ;
        RECT 2.97 1.5 3.445 1.56 ;
    END
    ANTENNAGATEAREA 0.675 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER li1 ;
  END A

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 4.125 6.17 4.385 ;
    END
  END vpb

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
    END
  END vpwr

  PIN lowlvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 6.17 2.945 ;
    END
  END lowlvpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 6.24 6.905 ;
    END
  END vgnd
  OBS
    LAYER li1 ;
      RECT 3.06 4.77 3.73 5.02 ;
      RECT 3.06 2.98 3.3 4.77 ;
      RECT 2.56 2.74 3.3 2.98 ;
      RECT 2.56 0.735 2.8 2.74 ;
      RECT 0 3.245 1.89 3.415 ;
      RECT 4.005 5.36 4.195 6.31 ;
      RECT 3.145 5.19 5.19 5.36 ;
      RECT 3.145 5.36 3.335 6.31 ;
      RECT 4.6 5.01 5.19 5.19 ;
      RECT 4.365 5.53 5.035 6.575 ;
      RECT 0 6.575 6.24 6.745 ;
      RECT 3.505 5.53 3.835 6.575 ;
      RECT 0.135 5.59 0.305 6.575 ;
      RECT 2.645 5.53 2.975 6.575 ;
      RECT 5.935 5.88 6.105 6.575 ;
      RECT 4.02 3.525 4.19 4.065 ;
      RECT 4.02 3.355 4.64 3.525 ;
      RECT 4.47 1.82 4.64 3.355 ;
      RECT 2.06 3.27 2.81 3.94 ;
      RECT 2.06 2.945 2.39 3.27 ;
      RECT 1.38 2.675 2.39 2.945 ;
      RECT 2.06 1.9 2.39 2.675 ;
      RECT 4.89 3.245 6.24 3.415 ;
      RECT 5.855 1.82 6.085 3.245 ;
      RECT 4.89 3.415 5.12 4.84 ;
      RECT 4.89 1.82 5.12 3.245 ;
      RECT 0 -0.085 6.24 0.085 ;
      RECT 5.76 0.085 6.09 1.13 ;
      RECT 3.115 0.085 3.445 1.13 ;
      RECT 3.975 0.085 4.305 1.05 ;
      RECT 4.835 0.085 5.165 1.13 ;
      RECT 2.02 0.085 2.35 1.13 ;
      RECT 0.135 0.085 0.305 1.07 ;
      RECT 3.68 3.185 3.85 4.235 ;
      RECT 3.615 1.22 4.665 1.39 ;
      RECT 3.615 0.35 3.805 1.22 ;
      RECT 4.475 0.35 4.665 1.22 ;
      RECT 4.39 4.405 4.72 4.84 ;
      RECT 3.68 4.235 4.72 4.405 ;
      RECT 4.39 3.695 4.72 4.235 ;
      RECT 4.02 1.39 4.19 3.015 ;
      RECT 3.68 3.015 4.19 3.185 ;
      RECT 0.1 3.65 0.33 4.4 ;
      RECT 5.91 3.65 6.14 4.4 ;
      RECT 5.205 5.72 5.55 6.31 ;
      RECT 5.205 5.53 5.865 5.72 ;
      RECT 5.36 5.05 5.865 5.53 ;
      RECT 5.36 3.68 5.55 5.05 ;
    LAYER mcon ;
      RECT 5.94 4.17 6.11 4.34 ;
      RECT 0.13 4.17 0.3 4.34 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 1.42 2.725 1.59 2.895 ;
      RECT 1.78 2.725 1.95 2.895 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 3.035 6.575 3.205 6.745 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.14 2.715 2.31 2.885 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
  END
END scs8ls_lpflow_lsbuf_lh_isowell_tap_2

MACRO scs8ls_lpflow_lsbuf_lh_isowell_tap_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.24 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.36 1.55 5.635 2.98 ;
        RECT 5.335 0.35 5.635 1.55 ;
    END
    ANTENNADIFFAREA 0.5041 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45 LAYER li1 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.83 3.29 2.15 ;
        RECT 2.97 1.56 3.63 1.83 ;
        RECT 2.97 1.5 3.445 1.56 ;
    END
  END A

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 4.125 6.17 4.385 ;
    END
  END vpb

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
    END
  END vpwr

  PIN lowlvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 6.17 2.945 ;
    END
  END lowlvpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 6.24 6.905 ;
    END
  END vgnd
  OBS
    LAYER li1 ;
      RECT 4.005 5.36 4.195 6.31 ;
      RECT 3.145 5.19 5.19 5.36 ;
      RECT 3.145 5.36 3.335 6.31 ;
      RECT 4.6 5.01 5.19 5.19 ;
      RECT 4.365 5.53 5.035 6.575 ;
      RECT 0 6.575 6.24 6.745 ;
      RECT 3.505 5.53 3.835 6.575 ;
      RECT 2.645 5.53 2.975 6.575 ;
      RECT 0.135 5.59 0.305 6.575 ;
      RECT 5.935 5.88 6.105 6.575 ;
      RECT 0.1 3.65 0.33 4.4 ;
      RECT 4.02 3.525 4.19 4.065 ;
      RECT 4.02 3.355 4.64 3.525 ;
      RECT 4.47 1.82 4.64 3.355 ;
      RECT 2.06 3.27 2.81 3.94 ;
      RECT 2.06 2.945 2.39 3.27 ;
      RECT 1.38 2.675 2.39 2.945 ;
      RECT 2.06 1.9 2.39 2.675 ;
      RECT 4.89 3.245 6.24 3.415 ;
      RECT 4.89 3.415 5.12 4.84 ;
      RECT 4.89 1.82 5.12 3.245 ;
      RECT 0 -0.085 6.24 0.085 ;
      RECT 5.935 0.085 6.105 1.07 ;
      RECT 3.115 0.085 3.445 1.13 ;
      RECT 3.975 0.085 4.305 1.05 ;
      RECT 4.835 0.085 5.165 1.13 ;
      RECT 0.135 0.085 0.305 1.07 ;
      RECT 2.02 0.085 2.35 1.13 ;
      RECT 5.91 3.65 6.14 4.4 ;
      RECT 3.68 3.185 3.85 4.235 ;
      RECT 3.615 1.22 4.665 1.39 ;
      RECT 3.615 0.35 3.805 1.22 ;
      RECT 4.475 0.35 4.665 1.22 ;
      RECT 4.39 4.405 4.72 4.84 ;
      RECT 3.68 4.235 4.72 4.405 ;
      RECT 4.39 3.695 4.72 4.235 ;
      RECT 4.02 1.39 4.19 3.015 ;
      RECT 3.68 3.015 4.19 3.185 ;
      RECT 5.205 5.72 5.55 6.31 ;
      RECT 5.205 5.53 5.865 5.72 ;
      RECT 5.36 5.05 5.865 5.53 ;
      RECT 5.36 3.68 5.55 5.05 ;
      RECT 3.06 4.77 3.73 5.02 ;
      RECT 3.06 2.98 3.3 4.77 ;
      RECT 2.56 2.74 3.3 2.98 ;
      RECT 2.56 0.735 2.8 2.74 ;
      RECT 0 3.245 1.89 3.415 ;
    LAYER mcon ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 0.13 4.17 0.3 4.34 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 1.42 2.725 1.59 2.895 ;
      RECT 1.78 2.725 1.95 2.895 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 3.035 6.575 3.205 6.745 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.14 2.715 2.31 2.885 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.94 4.17 6.11 4.34 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
  END
END scs8ls_lpflow_lsbuf_lh_isowell_tap_1

MACRO scs8ls_lpflow_srsdfxtp2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 15.36 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.47 4.305 1.795 ;
        RECT 4.025 1.125 4.305 1.47 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.134 LAYER li1 ;
  END SCD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.495 1.61 14.785 3.015 ;
        RECT 13.575 1.32 14.785 1.61 ;
        RECT 13.575 0.37 13.865 1.32 ;
        RECT 14.495 0.37 14.785 1.32 ;
        RECT 13.575 1.61 13.865 3.015 ;
    END
    ANTENNADIFFAREA 1.1088 ;
    ANTENNAPARTIALMETALSIDEAREA 1.174 LAYER li1 ;
  END Q

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045 5.035 1.69 5.455 ;
    END
    ANTENNAGATEAREA 0.318 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.145 LAYER li1 ;
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.095 0.455 1.765 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.84 5.205 5.17 5.875 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END CLK

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.86 5.205 7.45 5.445 ;
        RECT 6.23 5.445 7.45 5.535 ;
        RECT 6.23 5.535 7.015 5.615 ;
        RECT 6.23 5.615 6.4 6.235 ;
        RECT 3.72 6.235 6.4 6.405 ;
        RECT 3.72 5.455 3.95 6.235 ;
        RECT 3.59 5.225 3.95 5.455 ;
        RECT 3.59 4.8 3.92 5.225 ;
    END
    ANTENNAGATEAREA 0.598 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.231 LAYER li1 ;
  END SLEEPB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 15.36 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 15.36 6.905 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 15.36 3.575 ;
        RECT 9.295 2.985 9.945 3.085 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 3.715 15.29 3.985 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 10.715 6.575 10.885 6.745 ;
      RECT 14.235 3.27 14.405 3.44 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 6.575 10.405 6.745 ;
      RECT 14.595 3.245 14.765 3.415 ;
      RECT 10.1 3.785 10.27 3.955 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 9.755 6.575 9.925 6.745 ;
      RECT 9.74 3.785 9.91 3.955 ;
      RECT 9.715 3.03 9.885 3.2 ;
      RECT 9.355 3.03 9.525 3.2 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 6.575 9.445 6.745 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 6.575 8.965 6.745 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 6.575 8.485 6.745 ;
      RECT 8.175 3.245 8.345 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 6.575 8.005 6.745 ;
      RECT 7.815 3.18 7.985 3.35 ;
      RECT 7.455 3.18 7.625 3.35 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 6.575 14.725 6.745 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 6.575 7.525 6.745 ;
      RECT 7.095 3.18 7.265 3.35 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 6.575 7.045 6.745 ;
      RECT 6.825 3.765 6.995 3.935 ;
      RECT 6.735 3.18 6.905 3.35 ;
      RECT 6.465 3.765 6.635 3.935 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 6.575 6.565 6.745 ;
      RECT 6.375 3.18 6.545 3.35 ;
      RECT 6.015 3.18 6.185 3.35 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 13.115 6.575 13.285 6.745 ;
      RECT 5.155 3.745 5.325 3.915 ;
      RECT 12.795 3.27 12.965 3.44 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 4.795 3.785 4.965 3.955 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 4.115 3.115 4.285 3.285 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 3.755 3.115 3.925 3.285 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 13.875 3.27 14.045 3.44 ;
      RECT 3.395 3.115 3.565 3.285 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 13.515 3.27 13.685 3.44 ;
      RECT 3.035 3.115 3.205 3.285 ;
      RECT 3.035 6.575 3.205 6.745 ;
      RECT 13.595 6.575 13.765 6.745 ;
      RECT 2.675 3.115 2.845 3.285 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 13.155 3.27 13.325 3.44 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 2.315 3.115 2.485 3.285 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 14.075 6.575 14.245 6.745 ;
      RECT 1.955 3.245 2.125 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 6.575 12.805 6.745 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 15.035 6.575 15.205 6.745 ;
      RECT 15.075 3.245 15.245 3.415 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 12.155 6.575 12.325 6.745 ;
      RECT 11.9 3.345 12.07 3.515 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 6.575 11.845 6.745 ;
      RECT 11.54 3.345 11.71 3.515 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 6.575 11.365 6.745 ;
      RECT 10.715 -0.085 10.885 0.085 ;
    LAYER li1 ;
      RECT 8.3 6.19 9.9 6.39 ;
      RECT 9.73 5.55 9.9 6.19 ;
      RECT 9.73 5.38 10.87 5.55 ;
      RECT 10.7 5.55 10.87 6.19 ;
      RECT 9.945 5.285 10.275 5.38 ;
      RECT 10.7 6.19 12.025 6.39 ;
      RECT 11.695 5.865 12.025 6.19 ;
      RECT 11.695 5.525 12.005 5.865 ;
      RECT 6.06 5.035 6.69 5.275 ;
      RECT 6.57 3.985 6.9 4.695 ;
      RECT 6.465 3.705 7.005 3.985 ;
      RECT 6.04 3.795 6.295 4.155 ;
      RECT 6.04 4.155 6.35 4.605 ;
      RECT 5.72 4.605 6.35 4.775 ;
      RECT 5.72 4.775 5.89 5.475 ;
      RECT 5.38 5.475 5.89 5.69 ;
      RECT 5.38 5.69 6.06 6.065 ;
      RECT 10.55 3.755 10.88 4.94 ;
      RECT 9.36 4.94 12.05 5.11 ;
      RECT 9.36 5.11 9.61 5.24 ;
      RECT 11.05 5.11 11.3 6.02 ;
      RECT 9.36 4.91 9.61 4.94 ;
      RECT 11.72 5.11 12.05 5.19 ;
      RECT 11.72 4.875 12.05 4.94 ;
      RECT 9.02 3.775 9.395 4.685 ;
      RECT 9.02 3.605 9.475 3.775 ;
      RECT 9.02 4.685 9.19 5.69 ;
      RECT 9.305 3.585 9.475 3.605 ;
      RECT 9.02 5.69 9.36 6.02 ;
      RECT 9.305 3.415 11.22 3.585 ;
      RECT 11.05 3.585 11.22 3.635 ;
      RECT 11.05 3.635 11.33 4.305 ;
      RECT 9.305 2.985 9.935 3.245 ;
      RECT 9.41 1.885 9.74 2.985 ;
      RECT 10.02 3.985 10.35 4.685 ;
      RECT 9.69 3.755 10.35 3.985 ;
      RECT 12.585 4.985 14.555 5.155 ;
      RECT 14.225 5.155 14.555 6.05 ;
      RECT 12.585 3.87 12.825 4.985 ;
      RECT 12.28 3.67 12.825 3.87 ;
      RECT 12.28 2.635 12.59 3.67 ;
      RECT 12.585 5.155 12.755 5.33 ;
      RECT 12.175 5.33 12.755 5.5 ;
      RECT 12.175 5.5 12.425 5.685 ;
      RECT 14.05 4.275 14.38 4.985 ;
      RECT 12.76 3.415 14.5 3.465 ;
      RECT 12.76 3.245 15.36 3.415 ;
      RECT 14.955 1.855 15.245 3.245 ;
      RECT 13.2 3.5 13.53 4.605 ;
      RECT 12.76 3.465 13.53 3.5 ;
      RECT 12.76 2.25 13.405 3.245 ;
      RECT 12.415 1.92 13.405 2.25 ;
      RECT 12.75 1.855 13.405 1.92 ;
      RECT 14.035 1.855 14.325 3.245 ;
      RECT 11.725 3.57 12.11 4.4 ;
      RECT 11.5 3.305 12.11 3.57 ;
      RECT 0.155 5.255 0.805 5.955 ;
      RECT 0.595 4.17 0.805 5.255 ;
      RECT 0 -0.085 15.36 0.085 ;
      RECT 14.955 0.085 15.215 1.15 ;
      RECT 4.585 0.085 4.915 0.955 ;
      RECT 6.74 0.085 7.07 0.965 ;
      RECT 9.34 0.085 9.66 0.97 ;
      RECT 12.38 0.085 13.405 1.07 ;
      RECT 0.965 0.085 1.215 1.01 ;
      RECT 3.265 0.085 3.515 0.96 ;
      RECT 14.035 0.085 14.325 1.15 ;
      RECT 0 3.245 4.315 3.285 ;
      RECT 1.015 3.085 4.315 3.245 ;
      RECT 3.055 2.775 4.315 3.085 ;
      RECT 3.975 2.615 4.315 2.775 ;
      RECT 3.975 1.965 4.645 2.615 ;
      RECT 0 3.285 2.62 3.415 ;
      RECT 0.095 1.935 0.425 3.245 ;
      RECT 0.095 3.415 0.425 4.84 ;
      RECT 2.29 3.415 2.62 4.775 ;
      RECT 1.015 1.905 1.345 3.085 ;
      RECT 3.055 1.935 3.385 2.775 ;
      RECT 0 6.575 15.36 6.745 ;
      RECT 6.57 5.785 6.9 6.575 ;
      RECT 10.16 5.72 10.53 6.575 ;
      RECT 7.96 5.69 8.13 6.575 ;
      RECT 12.925 5.72 13.685 6.575 ;
      RECT 12.925 5.355 13.215 5.72 ;
      RECT 1.065 5.625 1.68 6.575 ;
      RECT 2.29 5.625 2.62 6.575 ;
      RECT 3.22 5.625 3.55 6.575 ;
      RECT 3.685 0.625 4.305 0.955 ;
      RECT 2.6 1.3 2.93 1.765 ;
      RECT 2.6 1.13 3.855 1.3 ;
      RECT 2.6 1.125 2.93 1.13 ;
      RECT 3.555 1.3 3.795 2.605 ;
      RECT 3.685 0.955 3.855 1.13 ;
      RECT 2.135 0.925 2.345 1.905 ;
      RECT 1.675 0.6 2.805 0.925 ;
      RECT 1.555 1.905 2.345 1.935 ;
      RECT 2.075 0.255 2.405 0.6 ;
      RECT 1.555 1.935 2.845 2.18 ;
      RECT 1.555 2.18 1.765 2.575 ;
      RECT 2.635 2.18 2.845 2.605 ;
      RECT 0.625 1.35 0.845 2.575 ;
      RECT 0.625 1.18 1.88 1.35 ;
      RECT 1.55 1.35 1.88 1.735 ;
      RECT 1.55 1.095 1.88 1.18 ;
      RECT 0.625 0.925 0.795 1.18 ;
      RECT 0.095 0.595 0.795 0.925 ;
      RECT 7.22 1.475 8.38 1.665 ;
      RECT 7.58 0.61 7.82 1.475 ;
      RECT 7.22 1.665 7.43 2.03 ;
      RECT 8.07 1.665 8.38 2.145 ;
      RECT 7.18 2.03 7.43 2.36 ;
      RECT 4.815 1.135 7.41 1.305 ;
      RECT 7.24 0.425 7.41 1.135 ;
      RECT 7.24 0.255 9.17 0.425 ;
      RECT 9 0.425 9.17 1.14 ;
      RECT 9 1.14 10 1.31 ;
      RECT 9.165 1.31 9.835 1.375 ;
      RECT 9.83 0.425 10 1.14 ;
      RECT 9.83 0.255 11.155 0.425 ;
      RECT 10.985 0.425 11.155 0.465 ;
      RECT 10.985 0.465 11.295 1.135 ;
      RECT 2.79 3.625 2.96 4.945 ;
      RECT 2.2 4.945 2.96 5.115 ;
      RECT 2.2 5.115 2.71 5.365 ;
      RECT 4.815 1.305 5.025 3.08 ;
      RECT 4.485 3.08 5.025 3.29 ;
      RECT 5.085 0.625 5.295 1.135 ;
      RECT 4.485 3.29 4.655 3.455 ;
      RECT 2.79 3.455 4.655 3.625 ;
      RECT 8.55 1.265 8.75 2.36 ;
      RECT 8.1 0.97 8.75 1.265 ;
      RECT 8.1 0.61 8.83 0.97 ;
      RECT 8.1 0.595 8.38 0.61 ;
      RECT 10.21 1.335 13.405 1.505 ;
      RECT 10.21 0.64 10.46 1.335 ;
      RECT 11.62 1.25 13.405 1.335 ;
      RECT 10.21 1.505 10.55 1.545 ;
      RECT 11.585 1.505 13.405 1.58 ;
      RECT 11.62 0.72 11.95 1.25 ;
      RECT 8.965 1.545 10.55 1.715 ;
      RECT 11.585 1.58 11.865 2.635 ;
      RECT 8.965 1.715 9.135 3.105 ;
      RECT 10.3 1.715 10.55 2.52 ;
      RECT 11.38 2.635 12.045 2.965 ;
      RECT 8.805 3.105 9.135 3.435 ;
      RECT 1.455 3.84 1.785 4.67 ;
      RECT 0.86 3.585 1.785 3.84 ;
      RECT 1.455 4.67 2.03 4.84 ;
      RECT 1.86 4.84 2.03 5.625 ;
      RECT 1.86 5.625 2.11 5.955 ;
      RECT 5.495 2.895 5.665 4.265 ;
      RECT 5.495 2.225 5.825 2.895 ;
      RECT 5.38 4.265 5.665 4.435 ;
      RECT 5.38 4.435 5.55 4.865 ;
      RECT 4.5 4.865 5.55 5.035 ;
      RECT 4.5 5.035 4.67 5.58 ;
      RECT 4.5 4.135 4.835 4.865 ;
      RECT 4.3 5.58 4.67 5.955 ;
      RECT 5.005 3.985 5.21 4.695 ;
      RECT 5.005 3.965 5.325 3.985 ;
      RECT 4.09 3.795 5.325 3.965 ;
      RECT 4.09 3.965 4.33 4.705 ;
      RECT 4.78 3.745 5.325 3.795 ;
      RECT 3.59 3.925 3.92 4.17 ;
      RECT 3.14 4.17 3.92 4.59 ;
      RECT 3.14 4.59 3.42 5.285 ;
      RECT 2.88 5.285 3.42 5.455 ;
      RECT 2.88 5.455 3.05 5.625 ;
      RECT 2.8 5.625 3.05 5.955 ;
      RECT 5.925 3.35 7.405 3.43 ;
      RECT 5.925 3.095 8.37 3.35 ;
      RECT 8.09 3.35 8.37 4.685 ;
      RECT 7.6 3.085 8.37 3.095 ;
      RECT 7.6 2.03 7.895 3.085 ;
      RECT 7.175 4.11 7.43 4.155 ;
      RECT 7.175 3.795 7.92 4.11 ;
      RECT 7.1 4.155 7.43 4.865 ;
      RECT 7.575 3.52 7.92 3.795 ;
      RECT 6.52 4.865 7.79 4.945 ;
      RECT 6.06 4.945 7.79 5.035 ;
      RECT 7.62 5.035 7.79 5.35 ;
      RECT 7.62 5.35 8.47 5.52 ;
      RECT 7.62 5.52 7.79 5.705 ;
      RECT 8.3 5.52 8.47 6.19 ;
      RECT 7.44 5.705 7.79 6.035 ;
  END
END scs8ls_lpflow_srsdfxtp2_4

MACRO scs8ls_lpflow_srsdfstp2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 17.28 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.32 1.145 5.625 1.815 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.059 LAYER li1 ;
  END SCD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.475 1.395 16.685 1.685 ;
        RECT 16.395 1.685 16.685 3.015 ;
        RECT 15.475 0.37 15.765 1.395 ;
        RECT 16.395 0.37 16.685 1.395 ;
        RECT 15.475 1.685 15.765 3.015 ;
    END
    ANTENNADIFFAREA 1.1088 ;
    ANTENNAPARTIALMETALSIDEAREA 1.174 LAYER li1 ;
  END Q

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.1 4.695 1.42 5.365 ;
    END
    ANTENNAGATEAREA 0.318 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.13 LAYER li1 ;
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.145 0.455 1.815 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.3 5.205 6.61 5.875 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.06 LAYER li1 ;
  END CLK

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.3 5.205 8.89 5.43 ;
        RECT 7.64 5.43 8.89 5.535 ;
        RECT 7.64 5.535 8.485 5.6 ;
        RECT 7.64 5.6 7.81 6.235 ;
        RECT 5.305 6.235 7.81 6.405 ;
        RECT 5.305 5.525 5.475 6.235 ;
        RECT 5.145 4.885 5.475 5.525 ;
    END
    ANTENNAGATEAREA 0.598 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.191 LAYER li1 ;
  END SLEEPB

  PIN SETB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met1 ;
        RECT 2.14 2.705 14.915 2.845 ;
        RECT 14.265 2.845 14.915 2.92 ;
        RECT 14.265 2.69 14.915 2.705 ;
        RECT 2.14 2.845 2.795 2.92 ;
        RECT 8.235 2.845 8.885 2.92 ;
        RECT 2.14 2.69 2.795 2.705 ;
        RECT 8.235 2.69 8.885 2.705 ;
    END
    ANTENNAGATEAREA 0.378 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 8.9915 LAYER met1 ;
  END SETB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 17.28 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 17.28 6.905 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 17.28 3.575 ;
        RECT 2.975 3.075 6.145 3.085 ;
        RECT 11.85 2.985 13.33 3.085 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 3.715 17.21 3.985 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 2.56 2.72 2.73 2.89 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 2.2 2.72 2.37 2.89 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.515 6.575 15.685 6.745 ;
      RECT 16.595 3.245 16.765 3.415 ;
      RECT 15.155 3.245 15.325 3.415 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 16.955 6.575 17.125 6.745 ;
      RECT 15.035 6.575 15.205 6.745 ;
      RECT 16.955 3.245 17.125 3.415 ;
      RECT 15.875 3.245 16.045 3.415 ;
      RECT 14.685 2.72 14.855 2.89 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 15.995 6.575 16.165 6.745 ;
      RECT 14.555 6.575 14.725 6.745 ;
      RECT 14.325 2.72 14.495 2.89 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 6.575 14.245 6.745 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 6.575 13.765 6.745 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 6.575 13.285 6.745 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 12.97 3.375 13.14 3.545 ;
      RECT 12.645 3.03 12.815 3.2 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 6.575 12.805 6.745 ;
      RECT 12.285 3.03 12.455 3.2 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 6.575 12.325 6.745 ;
      RECT 11.915 3.03 12.085 3.2 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 6.575 11.845 6.745 ;
      RECT 11.54 3.785 11.71 3.955 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 6.575 11.365 6.745 ;
      RECT 11.18 3.785 11.35 3.955 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 6.575 10.885 6.745 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 6.575 10.405 6.745 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 16.235 3.245 16.405 3.415 ;
      RECT 16.475 6.575 16.645 6.745 ;
      RECT 16.955 -0.085 17.125 0.085 ;
      RECT 9.755 6.575 9.925 6.745 ;
      RECT 9.615 3.245 9.785 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 6.575 9.445 6.745 ;
      RECT 9.255 3.18 9.425 3.35 ;
      RECT 8.895 3.18 9.065 3.35 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 6.575 8.965 6.745 ;
      RECT 8.655 2.72 8.825 2.89 ;
      RECT 8.535 3.18 8.705 3.35 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 6.575 8.485 6.745 ;
      RECT 8.295 2.72 8.465 2.89 ;
      RECT 8.255 3.765 8.425 3.935 ;
      RECT 8.175 3.18 8.345 3.35 ;
      RECT 7.895 3.765 8.065 3.935 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 6.575 8.005 6.745 ;
      RECT 7.815 3.18 7.985 3.35 ;
      RECT 7.455 3.18 7.625 3.35 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 7.355 6.575 7.525 6.745 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 6.575 7.045 6.745 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 6.575 6.565 6.745 ;
      RECT 6.155 3.785 6.325 3.955 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.105 6.085 3.275 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 5.555 3.105 5.725 3.275 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 5.265 3.785 5.435 3.955 ;
      RECT 5.195 3.105 5.365 3.275 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 4.835 3.105 5.005 3.275 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.105 4.645 3.275 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 4.115 3.105 4.285 3.275 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 3.755 3.105 3.925 3.275 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 3.395 3.105 3.565 3.275 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.105 3.205 3.275 ;
      RECT 3.035 6.575 3.205 6.745 ;
    LAYER li1 ;
      RECT 7.365 5.035 8.035 5.26 ;
      RECT 7.365 3.09 9.81 3.535 ;
      RECT 9.005 2.855 9.81 3.09 ;
      RECT 9.53 3.535 9.81 4.685 ;
      RECT 9.005 2.505 10.385 2.855 ;
      RECT 9.005 2.345 9.175 2.505 ;
      RECT 10.045 1.99 10.385 2.505 ;
      RECT 8.66 2.05 9.175 2.345 ;
      RECT 8.245 2.54 8.835 2.92 ;
      RECT 7.965 3.985 8.355 4.695 ;
      RECT 7.89 3.705 8.43 3.985 ;
      RECT 7.465 4.155 7.795 4.525 ;
      RECT 7.465 3.795 7.72 4.155 ;
      RECT 7.01 4.525 7.795 4.695 ;
      RECT 7.01 4.695 7.18 5.475 ;
      RECT 6.82 5.475 7.18 5.69 ;
      RECT 6.82 5.69 7.47 6.065 ;
      RECT 5.645 4.865 6.695 5.035 ;
      RECT 6.525 4.23 6.695 4.865 ;
      RECT 6.525 4.06 6.97 4.23 ;
      RECT 6.8 2.895 6.97 4.06 ;
      RECT 6.8 2.225 7.13 2.895 ;
      RECT 5.645 4.125 5.975 4.865 ;
      RECT 5.92 5.035 6.13 6.01 ;
      RECT 5.235 3.955 5.475 4.715 ;
      RECT 5.235 3.785 6.355 3.955 ;
      RECT 6.145 3.955 6.355 4.695 ;
      RECT 11.99 3.755 12.32 4.875 ;
      RECT 11.99 4.875 13.465 4.91 ;
      RECT 10.8 4.91 13.465 5.11 ;
      RECT 10.8 5.11 11.05 5.24 ;
      RECT 12.47 5.11 13.465 5.19 ;
      RECT 12.47 5.19 12.705 6.02 ;
      RECT 12.94 4.065 13.415 4.395 ;
      RECT 12.94 3.245 13.17 4.065 ;
      RECT 11.915 2.87 13.17 3.245 ;
      RECT 11.915 1.895 12.295 2.87 ;
      RECT 10.46 3.605 10.96 4.685 ;
      RECT 10.745 3.585 10.96 3.605 ;
      RECT 10.46 4.685 10.63 5.69 ;
      RECT 10.745 3.415 12.77 3.585 ;
      RECT 10.46 5.69 10.8 6.02 ;
      RECT 12.49 3.585 12.77 4.305 ;
      RECT 11.13 3.755 11.79 4.685 ;
      RECT 15.055 3.415 16.86 3.575 ;
      RECT 15.055 3.245 17.28 3.415 ;
      RECT 15.055 3.185 17.165 3.245 ;
      RECT 16.855 1.855 17.165 3.185 ;
      RECT 15.055 2.19 15.305 3.185 ;
      RECT 14.085 1.84 15.305 2.19 ;
      RECT 15.57 3.575 15.9 4.605 ;
      RECT 15.935 1.855 16.225 3.185 ;
      RECT 13.88 4.065 14.345 4.275 ;
      RECT 13.88 2.65 14.155 4.065 ;
      RECT 13.88 4.275 14.915 5.16 ;
      RECT 13.88 5.16 14.235 5.33 ;
      RECT 14.745 5.16 14.915 5.72 ;
      RECT 13.615 5.33 14.235 5.66 ;
      RECT 14.745 5.72 15.125 6.05 ;
      RECT 14.325 2.65 14.885 3.32 ;
      RECT 15.15 4.775 16.3 4.945 ;
      RECT 15.15 4.23 15.4 4.775 ;
      RECT 16.07 4.23 16.3 4.775 ;
      RECT 0 -0.085 17.28 0.085 ;
      RECT 16.855 0.085 17.105 1.15 ;
      RECT 5.88 0.085 6.21 0.955 ;
      RECT 9.21 0.085 10.115 0.86 ;
      RECT 11.99 0.085 15.305 0.285 ;
      RECT 11.99 0.285 12.645 0.94 ;
      RECT 14.045 0.285 15.305 1.125 ;
      RECT 0.965 0.085 1.3 1.06 ;
      RECT 2.93 0.085 3.25 1.015 ;
      RECT 4.56 0.085 4.81 0.975 ;
      RECT 15.935 0.085 16.225 1.15 ;
      RECT 6.38 0.255 8.73 0.425 ;
      RECT 8.56 0.425 8.73 1.03 ;
      RECT 8.56 1.03 10.455 1.125 ;
      RECT 7.925 1.125 10.455 1.2 ;
      RECT 10.285 0.425 10.455 1.03 ;
      RECT 7.925 1.2 8.73 1.295 ;
      RECT 10.285 0.255 11.82 0.425 ;
      RECT 7.925 1.295 8.515 1.455 ;
      RECT 11.65 0.425 11.82 1.11 ;
      RECT 11.65 1.11 13.09 1.345 ;
      RECT 12.835 1.345 13.09 2.31 ;
      RECT 3.85 3.615 4.02 4.945 ;
      RECT 2.825 4.945 4.02 5.115 ;
      RECT 2.825 5.115 3.335 5.365 ;
      RECT 6.38 0.425 6.63 3.445 ;
      RECT 3.85 3.445 6.63 3.615 ;
      RECT 0 6.575 17.28 6.745 ;
      RECT 8.01 6.265 9.57 6.575 ;
      RECT 11.51 5.72 11.96 6.575 ;
      RECT 14.28 6.22 16.315 6.575 ;
      RECT 8.01 5.77 8.6 6.265 ;
      RECT 9.4 5.72 9.57 6.265 ;
      RECT 14.28 5.83 14.575 6.22 ;
      RECT 15.985 5.72 16.315 6.22 ;
      RECT 14.405 5.33 14.575 5.83 ;
      RECT 1.1 6.28 4.11 6.575 ;
      RECT 4.73 5.68 5.06 6.575 ;
      RECT 2.05 5.625 2.315 6.28 ;
      RECT 2.915 5.625 3.245 6.28 ;
      RECT 3.845 5.625 4.11 6.28 ;
      RECT 1.1 5.605 1.395 6.28 ;
      RECT 0.625 1.615 1.8 1.82 ;
      RECT 0.625 0.975 0.795 1.615 ;
      RECT 1.55 1.145 1.8 1.615 ;
      RECT 0.625 1.82 0.845 2.66 ;
      RECT 0.095 0.645 0.795 0.975 ;
      RECT 1.97 0.975 2.19 1.99 ;
      RECT 1.675 0.255 2.325 0.975 ;
      RECT 1.515 1.99 2.19 2.175 ;
      RECT 1.515 2.175 1.785 2.66 ;
      RECT 4.98 0.645 5.6 0.975 ;
      RECT 3.975 1.32 4.225 1.815 ;
      RECT 3.975 1.145 5.15 1.32 ;
      RECT 4.85 1.32 5.1 2.655 ;
      RECT 4.98 0.975 5.15 1.145 ;
      RECT 3.585 0.975 3.805 1.985 ;
      RECT 3.45 0.255 4.1 0.975 ;
      RECT 3.585 1.985 4.14 2.205 ;
      RECT 3.91 2.205 4.14 2.655 ;
      RECT 2.495 1.185 3.415 1.855 ;
      RECT 2.495 0.65 2.76 1.185 ;
      RECT 2.495 1.855 2.76 2.34 ;
      RECT 7.575 1.185 7.755 1.71 ;
      RECT 7.305 0.955 7.755 1.185 ;
      RECT 7.575 1.71 9.615 1.88 ;
      RECT 7.305 0.595 8.39 0.955 ;
      RECT 8.28 1.88 8.49 2.345 ;
      RECT 9.345 1.88 9.615 2.335 ;
      RECT 11.145 1.515 12.665 1.725 ;
      RECT 11.145 0.595 11.48 1.515 ;
      RECT 11.145 1.725 11.46 3.025 ;
      RECT 12.465 1.725 12.665 2.48 ;
      RECT 10.225 3.025 11.46 3.245 ;
      RECT 12.465 2.48 13.67 2.7 ;
      RECT 10.225 3.245 10.575 3.435 ;
      RECT 13.26 1.625 13.67 2.48 ;
      RECT 13.34 2.7 13.67 3.68 ;
      RECT 13.26 1.295 15.305 1.625 ;
      RECT 13.26 0.755 13.565 1.295 ;
      RECT 10.585 1.59 10.895 2.38 ;
      RECT 10.045 1.54 10.895 1.59 ;
      RECT 9.065 1.37 10.895 1.54 ;
      RECT 10.625 0.625 10.895 1.37 ;
      RECT 0 3.245 1.345 3.415 ;
      RECT 0.095 2.84 1.345 3.245 ;
      RECT 1.015 1.99 1.345 2.84 ;
      RECT 0.16 3.415 0.52 4.84 ;
      RECT 0.095 2.02 0.455 2.84 ;
      RECT 0.69 4.17 0.93 5.255 ;
      RECT 0.235 5.255 0.93 5.955 ;
      RECT 2.895 3.275 3.265 4.775 ;
      RECT 2.895 3.24 6.21 3.275 ;
      RECT 2.93 2.855 6.21 3.24 ;
      RECT 2.93 2.025 3.28 2.855 ;
      RECT 4.315 2.835 6.21 2.855 ;
      RECT 4.315 1.985 4.68 2.835 ;
      RECT 5.27 2.015 6.21 2.835 ;
      RECT 4.215 3.925 4.995 4.595 ;
      RECT 4.215 4.595 4.54 5.285 ;
      RECT 3.505 5.285 4.54 5.455 ;
      RECT 3.505 5.455 3.675 5.535 ;
      RECT 4.28 5.455 4.54 5.955 ;
      RECT 3.415 5.535 3.675 5.955 ;
      RECT 2.14 2.61 2.76 2.94 ;
      RECT 1.59 3.84 1.99 4.64 ;
      RECT 0.895 3.585 1.99 3.84 ;
      RECT 1.59 4.64 2.655 4.84 ;
      RECT 1.59 4.84 1.88 5.955 ;
      RECT 2.485 4.84 2.655 5.535 ;
      RECT 2.485 5.535 2.745 5.955 ;
      RECT 8.525 4.155 9.36 4.865 ;
      RECT 8.6 3.795 9.36 4.155 ;
      RECT 7.365 4.865 9.36 5.035 ;
      RECT 9.03 3.73 9.36 3.795 ;
      RECT 9.06 5.035 9.36 5.38 ;
      RECT 9.06 5.38 9.91 5.55 ;
      RECT 9.06 5.55 9.23 5.705 ;
      RECT 9.74 5.55 9.91 6.19 ;
      RECT 8.77 5.705 9.23 6.065 ;
      RECT 9.74 6.19 11.34 6.39 ;
      RECT 11.17 5.55 11.34 6.19 ;
      RECT 11.17 5.38 12.3 5.55 ;
      RECT 12.13 5.55 12.3 6.19 ;
      RECT 11.225 5.285 12.3 5.38 ;
      RECT 12.13 6.19 13.445 6.39 ;
      RECT 13.135 5.525 13.445 6.19 ;
  END
END scs8ls_lpflow_srsdfstp2_4

MACRO scs8ls_lpflow_srsdfrtp2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 17.76 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.5 1.125 6.085 1.44 ;
        RECT 5.5 1.44 5.725 1.795 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.183 LAYER li1 ;
  END SCD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.895 1.615 17.185 3.015 ;
        RECT 16.055 1.345 17.185 1.615 ;
        RECT 16.055 1.615 16.325 1.82 ;
        RECT 16.055 0.37 16.325 1.345 ;
        RECT 16.895 0.37 17.185 1.345 ;
        RECT 15.975 1.82 16.325 2.09 ;
        RECT 15.975 2.09 16.255 3.015 ;
    END
    ANTENNADIFFAREA 1.1088 ;
    ANTENNAPARTIALMETALSIDEAREA 1.178 LAYER li1 ;
  END Q

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.49 5.035 2.08 5.455 ;
    END
    ANTENNAGATEAREA 0.318 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.134 LAYER li1 ;
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.095 0.425 1.765 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.058 LAYER li1 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.68 4.895 7.195 5.515 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.091 LAYER li1 ;
  END CLK

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.15 5.205 9.85 5.38 ;
        RECT 8.615 5.38 9.85 5.535 ;
        RECT 8.615 5.535 9.32 5.55 ;
        RECT 8.615 5.55 8.785 6.235 ;
        RECT 7.225 6.235 8.785 6.405 ;
        RECT 7.225 6.205 7.595 6.235 ;
        RECT 7.425 5.265 7.595 6.205 ;
        RECT 7.425 4.935 7.74 5.265 ;
    END
    ANTENNAGATEAREA 0.598 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.986 LAYER li1 ;
  END SLEEPB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 17.76 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 17.76 6.905 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 17.76 3.575 ;
        RECT 6.38 2.985 8.11 3.085 ;
        RECT 10.405 2.985 13.82 3.085 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 3.715 17.69 3.985 ;
    END
  END kapwr

  PIN RESETB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met1 ;
        RECT 2.535 2.705 15.33 2.845 ;
        RECT 14.67 2.845 15.33 2.935 ;
        RECT 15.015 2.69 15.33 2.705 ;
        RECT 2.535 2.845 3.215 2.935 ;
        RECT 8.45 2.845 9.1 2.92 ;
        RECT 2.535 2.69 3.215 2.705 ;
        RECT 8.45 2.69 9.1 2.705 ;
    END
    ANTENNAGATEAREA 0.378 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 9.0265 LAYER met1 ;
  END RESETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 13.23 3.065 13.4 3.235 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 6.575 13.285 6.745 ;
      RECT 12.87 3.015 13.04 3.185 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 6.575 12.805 6.745 ;
      RECT 12.51 3.015 12.68 3.185 ;
      RECT 12.5 3.785 12.67 3.955 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 6.575 12.325 6.745 ;
      RECT 12.14 3.785 12.31 3.955 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 6.575 11.845 6.745 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 6.575 11.365 6.745 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 6.575 10.885 6.745 ;
      RECT 10.51 3.375 10.68 3.545 ;
      RECT 10.465 3.015 10.635 3.185 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 6.575 10.405 6.745 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 6.575 9.925 6.745 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 6.575 9.445 6.745 ;
      RECT 9.215 3.765 9.385 3.935 ;
      RECT 8.87 2.72 9.04 2.89 ;
      RECT 8.855 3.765 9.025 3.935 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 6.575 8.965 6.745 ;
      RECT 8.51 2.72 8.68 2.89 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 6.575 8.485 6.745 ;
      RECT 8.04 3.785 8.21 3.955 ;
      RECT 7.88 3.105 8.05 3.275 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 6.575 8.005 6.745 ;
      RECT 7.68 3.785 7.85 3.955 ;
      RECT 7.52 3.105 7.69 3.275 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 6.575 7.525 6.745 ;
      RECT 7.16 3.105 7.33 3.275 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 6.575 7.045 6.745 ;
      RECT 6.8 3.105 6.97 3.275 ;
      RECT 6.795 3.785 6.965 3.955 ;
      RECT 6.44 3.015 6.61 3.185 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 6.575 6.565 6.745 ;
      RECT 6.315 3.375 6.485 3.545 ;
      RECT 15.635 3.295 15.805 3.465 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 17.435 3.245 17.605 3.415 ;
      RECT 5.475 3.245 5.645 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 5.105 3.245 5.275 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 4.525 3.245 4.695 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 4.155 3.245 4.325 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 3.785 3.245 3.955 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 17.435 -0.085 17.605 0.085 ;
      RECT 17.075 3.245 17.245 3.415 ;
      RECT 16.955 -0.085 17.125 0.085 ;
      RECT 16.955 6.575 17.125 6.745 ;
      RECT 17.435 6.575 17.605 6.745 ;
      RECT 16.715 3.245 16.885 3.415 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 16.475 6.575 16.645 6.745 ;
      RECT 16.355 3.295 16.525 3.465 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 6.575 16.165 6.745 ;
      RECT 15.995 3.295 16.165 3.465 ;
      RECT 15.1 2.735 15.27 2.905 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 6.575 15.685 6.745 ;
      RECT 14.74 2.735 14.91 2.905 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 6.575 15.205 6.745 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 6.575 14.725 6.745 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 3.415 3.245 3.585 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 6.575 3.205 6.745 ;
      RECT 2.985 2.735 3.155 2.905 ;
      RECT 2.595 2.735 2.765 2.905 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 1.26 3.245 1.43 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 0.89 3.245 1.06 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 0.525 3.245 0.695 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 14.075 6.575 14.245 6.745 ;
      RECT 13.95 3.375 14.12 3.545 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 6.575 13.765 6.745 ;
      RECT 13.59 3.065 13.76 3.235 ;
    LAYER li1 ;
      RECT 3.505 3.415 3.835 4.775 ;
      RECT 3.355 2.79 5.725 3.415 ;
      RECT 3.355 2.525 3.825 2.79 ;
      RECT 5.385 1.97 5.725 2.79 ;
      RECT 4.475 1.935 4.805 2.79 ;
      RECT 3.115 2.315 3.825 2.525 ;
      RECT 3.115 1.925 3.445 2.315 ;
      RECT 4.77 4.17 5.54 4.595 ;
      RECT 5.21 3.925 5.54 4.17 ;
      RECT 4.77 4.595 5.09 5.43 ;
      RECT 4.005 5.43 5.13 5.6 ;
      RECT 4.005 5.6 4.195 5.995 ;
      RECT 4.88 5.6 5.13 5.955 ;
      RECT 6.275 3.275 6.525 4.385 ;
      RECT 6.275 3.085 8.15 3.275 ;
      RECT 6.275 1.95 6.69 3.085 ;
      RECT 7.855 1.93 8.15 3.085 ;
      RECT 6.715 3.705 7.045 4.385 ;
      RECT 9.485 4.155 9.815 4.865 ;
      RECT 9.56 4.11 9.815 4.155 ;
      RECT 8.81 4.865 10.19 4.955 ;
      RECT 9.56 3.795 10.32 4.11 ;
      RECT 8.31 4.955 10.19 5.035 ;
      RECT 9.99 3.52 10.32 3.795 ;
      RECT 10.02 5.035 10.19 5.38 ;
      RECT 10.02 5.38 11.22 5.55 ;
      RECT 10.02 5.55 10.19 5.735 ;
      RECT 11.05 5.55 11.22 6.22 ;
      RECT 9.825 5.735 10.19 6.065 ;
      RECT 11.05 6.22 12.3 6.39 ;
      RECT 12.13 5.55 12.3 6.22 ;
      RECT 12.13 5.38 13.26 5.55 ;
      RECT 13.09 5.55 13.26 6.22 ;
      RECT 12.345 5.285 12.675 5.38 ;
      RECT 13.09 6.22 14.425 6.39 ;
      RECT 14.095 5.865 14.425 6.22 ;
      RECT 14.095 5.525 14.405 5.865 ;
      RECT 8.31 5.035 8.98 5.21 ;
      RECT 8.955 3.985 9.285 4.695 ;
      RECT 8.85 3.705 9.39 3.985 ;
      RECT 8.41 2.655 9.14 2.93 ;
      RECT 8.41 1.935 9.08 2.655 ;
      RECT 8.425 4.155 8.755 4.615 ;
      RECT 8.425 3.795 8.68 4.155 ;
      RECT 7.97 4.615 8.755 4.695 ;
      RECT 7.97 4.695 8.595 4.785 ;
      RECT 7.97 4.785 8.14 5.475 ;
      RECT 7.765 5.475 8.14 5.735 ;
      RECT 7.765 5.735 8.445 6.065 ;
      RECT 7.635 3.785 8.255 4.445 ;
      RECT 15.025 4.995 16.955 5.165 ;
      RECT 16.625 5.165 16.955 6.05 ;
      RECT 13.555 2.715 14.51 2.885 ;
      RECT 14.34 2.885 14.51 3.825 ;
      RECT 14.34 3.825 15.265 3.995 ;
      RECT 15.025 3.995 15.265 4.995 ;
      RECT 15.025 5.165 15.195 5.33 ;
      RECT 14.575 5.33 15.195 5.5 ;
      RECT 14.575 5.5 14.825 5.685 ;
      RECT 16.45 4.275 16.78 4.995 ;
      RECT 12.95 3.755 13.28 4.94 ;
      RECT 11.76 4.94 14.855 5.11 ;
      RECT 11.76 5.11 12.01 5.24 ;
      RECT 13.45 5.11 13.7 6.05 ;
      RECT 11.76 4.91 12.01 4.94 ;
      RECT 14.265 5.11 14.855 5.16 ;
      RECT 14.265 4.83 14.855 4.94 ;
      RECT 15.495 3.185 17.625 3.245 ;
      RECT 15.495 3.245 17.76 3.415 ;
      RECT 17.355 1.855 17.625 3.185 ;
      RECT 12.45 3.055 14.17 3.245 ;
      RECT 12.45 2.955 13.385 3.055 ;
      RECT 13.9 3.245 14.17 4.165 ;
      RECT 12.45 2.545 13.03 2.955 ;
      RECT 13.9 4.165 14.455 4.445 ;
      RECT 12.45 2.535 14.51 2.545 ;
      RECT 12.45 2.365 15.805 2.535 ;
      RECT 12.45 2.34 14.43 2.365 ;
      RECT 15.495 2.535 15.805 3.185 ;
      RECT 15.495 1.855 15.805 2.365 ;
      RECT 12.45 1.945 13.03 2.34 ;
      RECT 14.1 1.92 14.43 2.34 ;
      RECT 12.745 1.825 13.03 1.945 ;
      RECT 15.495 4.075 15.93 4.605 ;
      RECT 16.435 2.26 16.725 3.185 ;
      RECT 15.495 3.415 16.75 4.075 ;
      RECT 16.495 1.855 16.725 2.26 ;
      RECT 11.42 3.585 11.795 4.685 ;
      RECT 11.42 3.415 13.73 3.585 ;
      RECT 11.42 4.685 11.59 5.72 ;
      RECT 13.45 3.585 13.73 4.305 ;
      RECT 11.42 5.72 11.76 6.05 ;
      RECT 12.42 3.985 12.75 4.685 ;
      RECT 12.09 3.755 12.75 3.985 ;
      RECT 10.49 3.4 10.78 4.685 ;
      RECT 10.49 3.35 10.695 3.4 ;
      RECT 10.405 2.73 10.695 3.35 ;
      RECT 10.405 1.97 10.77 2.73 ;
      RECT 14.68 2.935 14.93 3.4 ;
      RECT 14.68 2.705 15.325 2.935 ;
      RECT 0 6.575 17.76 6.745 ;
      RECT 8.955 5.72 9.285 6.575 ;
      RECT 10.36 5.72 10.75 6.575 ;
      RECT 12.5 5.72 12.89 6.575 ;
      RECT 15.365 5.72 16.085 6.575 ;
      RECT 15.365 5.355 15.615 5.72 ;
      RECT 1.51 5.625 1.775 6.575 ;
      RECT 2.64 5.77 2.97 6.575 ;
      RECT 4.37 5.77 4.7 6.575 ;
      RECT 5.84 5.67 6.17 6.575 ;
      RECT 3.505 5.625 3.835 6.575 ;
      RECT 0 -0.085 17.76 0.085 ;
      RECT 17.355 0.085 17.655 1.15 ;
      RECT 6.02 0.085 6.35 0.86 ;
      RECT 8.115 0.085 8.325 0.94 ;
      RECT 10.415 0.085 11.825 0.97 ;
      RECT 14.67 0.085 14.92 0.81 ;
      RECT 15.585 0.085 15.885 1.15 ;
      RECT 1.03 0.085 1.36 0.97 ;
      RECT 3.085 0.085 3.405 0.99 ;
      RECT 4.615 0.085 4.935 1 ;
      RECT 16.495 0.085 16.725 1.15 ;
      RECT 2.115 0.925 2.325 1.935 ;
      RECT 2.115 0.895 2.39 0.925 ;
      RECT 1.62 1.935 2.325 2.145 ;
      RECT 1.74 0.57 2.39 0.895 ;
      RECT 1.62 2.145 1.91 2.605 ;
      RECT 2.14 0.255 2.39 0.57 ;
      RECT 0.69 1.35 0.91 2.605 ;
      RECT 0.69 1.18 1.945 1.35 ;
      RECT 1.615 1.35 1.945 1.735 ;
      RECT 1.615 1.125 1.945 1.18 ;
      RECT 0.69 0.925 0.86 1.18 ;
      RECT 0.16 0.595 0.86 0.925 ;
      RECT 2.495 1.095 2.915 1.825 ;
      RECT 2.645 0.64 2.915 1.095 ;
      RECT 2.66 1.825 2.915 2.34 ;
      RECT 5.105 0.625 5.805 0.955 ;
      RECT 4.02 1.63 4.35 1.735 ;
      RECT 4.02 1.415 5.33 1.63 ;
      RECT 4.975 1.63 5.215 2.605 ;
      RECT 4.02 1.125 4.35 1.415 ;
      RECT 5.105 0.955 5.33 1.415 ;
      RECT 3.64 0.925 3.85 1.935 ;
      RECT 3.575 0.6 4.225 0.925 ;
      RECT 3.64 1.935 4.265 2.145 ;
      RECT 3.575 0.255 3.825 0.6 ;
      RECT 4.055 2.145 4.265 2.605 ;
      RECT 8.495 0.255 10.245 0.425 ;
      RECT 10.075 0.425 10.245 1.15 ;
      RECT 10.075 1.15 12.165 1.32 ;
      RECT 10.075 1.32 10.925 1.46 ;
      RECT 11.995 0.425 12.165 1.15 ;
      RECT 11.995 0.255 13.18 0.425 ;
      RECT 13.01 0.425 13.18 0.465 ;
      RECT 13.01 0.465 13.28 1.135 ;
      RECT 5.895 1.61 6.69 1.78 ;
      RECT 6.52 0.425 6.69 1.61 ;
      RECT 5.895 1.78 6.105 3.585 ;
      RECT 4.035 3.585 6.105 3.755 ;
      RECT 5.775 3.755 6.105 4.155 ;
      RECT 5.71 4.155 6.105 4.365 ;
      RECT 5.71 4.365 5.92 5.29 ;
      RECT 5.46 5.29 5.92 5.5 ;
      RECT 5.46 5.5 5.67 6.02 ;
      RECT 4.035 3.755 4.205 4.945 ;
      RECT 3.335 4.945 4.205 5.115 ;
      RECT 3.335 5.115 4.005 5.26 ;
      RECT 6.52 0.255 7.945 0.425 ;
      RECT 7.775 0.425 7.945 1.12 ;
      RECT 7.775 1.12 8.665 1.29 ;
      RECT 8.495 0.425 8.665 1.12 ;
      RECT 9.98 1.63 11.22 1.8 ;
      RECT 9.98 1.8 10.15 3.135 ;
      RECT 10.94 1.8 11.22 2.69 ;
      RECT 8.51 3.135 10.15 3.305 ;
      RECT 6.34 5.685 7.255 6.015 ;
      RECT 6.18 4.725 6.51 5.21 ;
      RECT 6.34 5.21 6.51 5.685 ;
      RECT 7.295 3.615 7.465 3.705 ;
      RECT 7.215 3.705 7.465 4.555 ;
      RECT 6.18 4.555 7.465 4.725 ;
      RECT 8.51 3.305 8.68 3.445 ;
      RECT 7.295 3.445 8.68 3.615 ;
      RECT 9.38 1.305 9.55 1.93 ;
      RECT 9.19 0.94 9.55 1.305 ;
      RECT 9.25 1.93 9.55 2.26 ;
      RECT 8.835 0.595 9.905 0.94 ;
      RECT 7.395 1.665 7.655 2.26 ;
      RECT 7.395 1.475 9.21 1.665 ;
      RECT 8.54 1.665 9.21 1.725 ;
      RECT 7.395 0.61 7.605 1.475 ;
      RECT 6.86 0.61 7.1 2.645 ;
      RECT 6.86 2.645 7.685 2.895 ;
      RECT 13.25 1.65 13.58 2.17 ;
      RECT 13.25 1.48 15.885 1.65 ;
      RECT 13.25 1.475 13.7 1.48 ;
      RECT 14.95 1.65 15.28 2.195 ;
      RECT 15.295 1.32 15.885 1.48 ;
      RECT 12.335 1.305 13.7 1.475 ;
      RECT 12.335 1.475 12.575 1.49 ;
      RECT 12.335 0.625 12.575 1.305 ;
      RECT 13.45 0.48 13.7 1.305 ;
      RECT 11.85 1.49 12.575 1.775 ;
      RECT 11.85 1.775 12.18 2.9 ;
      RECT 10.865 2.9 12.18 3.07 ;
      RECT 10.865 3.07 11.455 3.23 ;
      RECT 14.2 0.98 15.35 1.15 ;
      RECT 14.2 0.48 14.5 0.98 ;
      RECT 15.09 0.48 15.35 0.98 ;
      RECT 0.925 3.585 2.61 3.84 ;
      RECT 2.25 3.84 2.61 4.845 ;
      RECT 2.25 4.845 2.46 5.43 ;
      RECT 2.25 5.43 3.335 5.6 ;
      RECT 2.25 5.6 2.46 5.955 ;
      RECT 3.145 5.6 3.335 5.995 ;
      RECT 0.505 4.11 0.87 4.84 ;
      RECT 0.505 3.415 0.725 4.11 ;
      RECT 0 3.245 1.46 3.415 ;
      RECT 0.22 2.79 1.46 3.245 ;
      RECT 0.22 2.785 1.41 2.79 ;
      RECT 0.22 1.935 0.5 2.785 ;
      RECT 1.08 1.935 1.41 2.785 ;
      RECT 1.08 4.17 1.32 5.255 ;
      RECT 0.6 5.255 1.32 5.925 ;
      RECT 1.08 5.925 1.32 5.955 ;
      RECT 2.565 2.695 3.185 3.025 ;
  END
END scs8ls_lpflow_srsdfrtp2_4

MACRO scs8ls_lpflow_srsdfxtp2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 14.88 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.47 4.305 1.795 ;
        RECT 4.025 1.125 4.305 1.47 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.134 LAYER li1 ;
  END SCD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.555 0.37 13.845 3.015 ;
    END
    ANTENNADIFFAREA 0.5544 ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1 ;
  END Q

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045 5.035 1.69 5.455 ;
    END
    ANTENNAGATEAREA 0.318 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.145 LAYER li1 ;
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.095 0.455 1.765 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.84 5.205 5.17 5.875 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END CLK

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.86 5.205 7.45 5.445 ;
        RECT 6.23 5.445 7.45 5.535 ;
        RECT 6.23 5.535 7.015 5.615 ;
        RECT 6.23 5.615 6.4 6.235 ;
        RECT 3.72 6.235 6.4 6.405 ;
        RECT 3.72 5.455 3.95 6.235 ;
        RECT 3.59 5.225 3.95 5.455 ;
        RECT 3.59 4.8 3.92 5.225 ;
    END
    ANTENNAGATEAREA 0.598 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.231 LAYER li1 ;
  END SLEEPB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.88 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 14.88 6.905 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.88 3.575 ;
        RECT 9.295 2.985 9.945 3.085 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 3.715 14.81 3.985 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 9.74 3.785 9.91 3.955 ;
      RECT 9.715 3.03 9.885 3.2 ;
      RECT 9.355 3.03 9.525 3.2 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 6.575 9.445 6.745 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 6.575 8.965 6.745 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 6.575 8.485 6.745 ;
      RECT 8.175 3.245 8.345 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 6.575 8.005 6.745 ;
      RECT 7.815 3.18 7.985 3.35 ;
      RECT 7.455 3.18 7.625 3.35 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 6.575 14.725 6.745 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 6.575 7.525 6.745 ;
      RECT 7.095 3.18 7.265 3.35 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 6.575 7.045 6.745 ;
      RECT 6.825 3.765 6.995 3.935 ;
      RECT 6.735 3.18 6.905 3.35 ;
      RECT 6.465 3.765 6.635 3.935 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 6.575 6.565 6.745 ;
      RECT 6.375 3.18 6.545 3.35 ;
      RECT 6.015 3.18 6.185 3.35 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 13.115 6.575 13.285 6.745 ;
      RECT 5.155 3.745 5.325 3.915 ;
      RECT 12.795 3.27 12.965 3.44 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 4.795 3.785 4.965 3.955 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 4.115 3.115 4.285 3.285 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 3.755 3.115 3.925 3.285 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 13.875 3.27 14.045 3.44 ;
      RECT 3.395 3.115 3.565 3.285 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 13.515 3.27 13.685 3.44 ;
      RECT 3.035 3.115 3.205 3.285 ;
      RECT 3.035 6.575 3.205 6.745 ;
      RECT 13.595 6.575 13.765 6.745 ;
      RECT 2.675 3.115 2.845 3.285 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 13.155 3.27 13.325 3.44 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 2.315 3.115 2.485 3.285 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 14.075 6.575 14.245 6.745 ;
      RECT 1.955 3.245 2.125 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 6.575 12.805 6.745 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 6.575 12.325 6.745 ;
      RECT 11.9 3.345 12.07 3.515 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 6.575 11.845 6.745 ;
      RECT 11.54 3.345 11.71 3.515 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 6.575 11.365 6.745 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 6.575 10.885 6.745 ;
      RECT 14.235 3.27 14.405 3.44 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 6.575 10.405 6.745 ;
      RECT 14.595 3.245 14.765 3.415 ;
      RECT 10.1 3.785 10.27 3.955 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 9.755 6.575 9.925 6.745 ;
    LAYER li1 ;
      RECT 11.05 5.11 11.3 6.02 ;
      RECT 11.72 5.11 12.05 5.19 ;
      RECT 11.72 4.875 12.05 4.94 ;
      RECT 9.02 3.775 9.395 4.685 ;
      RECT 9.02 3.605 9.475 3.775 ;
      RECT 9.02 4.685 9.19 5.69 ;
      RECT 9.305 3.585 9.475 3.605 ;
      RECT 9.02 5.69 9.36 6.02 ;
      RECT 9.305 3.415 11.22 3.585 ;
      RECT 11.05 3.585 11.22 3.635 ;
      RECT 11.05 3.635 11.33 4.305 ;
      RECT 9.305 2.985 9.935 3.245 ;
      RECT 9.41 1.885 9.74 2.985 ;
      RECT 7.175 4.11 7.43 4.155 ;
      RECT 7.175 3.795 7.92 4.11 ;
      RECT 7.1 4.155 7.43 4.865 ;
      RECT 7.575 3.52 7.92 3.795 ;
      RECT 6.52 4.865 7.79 4.945 ;
      RECT 6.06 4.945 7.79 5.035 ;
      RECT 7.62 5.035 7.79 5.35 ;
      RECT 7.62 5.35 8.47 5.52 ;
      RECT 7.62 5.52 7.79 5.705 ;
      RECT 8.3 5.52 8.47 6.19 ;
      RECT 7.44 5.705 7.79 6.035 ;
      RECT 8.3 6.19 9.9 6.39 ;
      RECT 9.73 5.55 9.9 6.19 ;
      RECT 9.73 5.38 10.87 5.55 ;
      RECT 10.7 5.55 10.87 6.19 ;
      RECT 9.945 5.285 10.275 5.38 ;
      RECT 10.7 6.19 12.025 6.39 ;
      RECT 11.695 5.865 12.025 6.19 ;
      RECT 11.695 5.525 12.005 5.865 ;
      RECT 6.06 5.035 6.69 5.275 ;
      RECT 10.02 3.985 10.35 4.685 ;
      RECT 9.69 3.755 10.35 3.985 ;
      RECT 12.76 3.415 14.5 3.465 ;
      RECT 12.76 3.245 14.88 3.415 ;
      RECT 14.015 1.855 14.305 3.245 ;
      RECT 13.2 3.5 13.53 4.605 ;
      RECT 12.76 3.465 13.53 3.5 ;
      RECT 12.76 2.25 13.345 3.245 ;
      RECT 12.415 1.92 13.345 2.25 ;
      RECT 13.095 1.855 13.345 1.92 ;
      RECT 11.725 3.57 12.11 4.4 ;
      RECT 11.5 3.305 12.11 3.57 ;
      RECT 12.585 4.985 14.555 5.155 ;
      RECT 14.225 5.155 14.555 6.05 ;
      RECT 14.05 4.275 14.38 4.985 ;
      RECT 12.585 3.87 12.825 4.985 ;
      RECT 12.28 3.67 12.825 3.87 ;
      RECT 12.28 2.635 12.59 3.67 ;
      RECT 12.585 5.155 12.755 5.33 ;
      RECT 12.175 5.33 12.755 5.5 ;
      RECT 12.175 5.5 12.425 5.685 ;
      RECT 0.155 5.255 0.805 5.955 ;
      RECT 0.595 4.17 0.805 5.255 ;
      RECT 0 -0.085 14.88 0.085 ;
      RECT 14.015 0.085 14.275 1.15 ;
      RECT 4.585 0.085 4.915 0.955 ;
      RECT 6.74 0.085 7.07 0.965 ;
      RECT 9.34 0.085 9.66 0.97 ;
      RECT 12.38 0.085 13.385 1.07 ;
      RECT 0.965 0.085 1.215 1.01 ;
      RECT 3.265 0.085 3.515 0.96 ;
      RECT 0 3.245 4.315 3.285 ;
      RECT 1.015 3.085 4.315 3.245 ;
      RECT 3.055 2.775 4.315 3.085 ;
      RECT 3.975 2.615 4.315 2.775 ;
      RECT 3.975 1.965 4.645 2.615 ;
      RECT 0 3.285 2.62 3.415 ;
      RECT 0.095 1.935 0.425 3.245 ;
      RECT 0.095 3.415 0.425 4.84 ;
      RECT 2.29 3.415 2.62 4.775 ;
      RECT 1.015 1.905 1.345 3.085 ;
      RECT 3.055 1.935 3.385 2.775 ;
      RECT 0 6.575 14.88 6.745 ;
      RECT 6.57 5.785 6.9 6.575 ;
      RECT 10.16 5.72 10.53 6.575 ;
      RECT 7.96 5.69 8.13 6.575 ;
      RECT 12.925 5.72 13.685 6.575 ;
      RECT 12.925 5.355 13.215 5.72 ;
      RECT 1.065 5.625 1.68 6.575 ;
      RECT 2.29 5.625 2.62 6.575 ;
      RECT 3.22 5.625 3.55 6.575 ;
      RECT 3.685 0.625 4.305 0.955 ;
      RECT 2.6 1.3 2.93 1.765 ;
      RECT 2.6 1.13 3.855 1.3 ;
      RECT 2.6 1.125 2.93 1.13 ;
      RECT 3.555 1.3 3.795 2.605 ;
      RECT 3.685 0.955 3.855 1.13 ;
      RECT 2.135 0.925 2.345 1.905 ;
      RECT 1.675 0.6 2.805 0.925 ;
      RECT 1.555 1.905 2.345 1.935 ;
      RECT 2.075 0.255 2.405 0.6 ;
      RECT 1.555 1.935 2.845 2.18 ;
      RECT 1.555 2.18 1.765 2.575 ;
      RECT 2.635 2.18 2.845 2.605 ;
      RECT 0.625 1.35 0.845 2.575 ;
      RECT 0.625 1.18 1.88 1.35 ;
      RECT 1.55 1.35 1.88 1.735 ;
      RECT 1.55 1.095 1.88 1.18 ;
      RECT 0.625 0.925 0.795 1.18 ;
      RECT 0.095 0.595 0.795 0.925 ;
      RECT 4.815 1.135 7.41 1.305 ;
      RECT 7.24 0.425 7.41 1.135 ;
      RECT 7.24 0.255 9.17 0.425 ;
      RECT 9 0.425 9.17 1.14 ;
      RECT 9 1.14 10 1.31 ;
      RECT 9.165 1.31 9.835 1.375 ;
      RECT 9.83 0.425 10 1.14 ;
      RECT 9.83 0.255 11.155 0.425 ;
      RECT 10.985 0.425 11.155 0.465 ;
      RECT 10.985 0.465 11.295 1.135 ;
      RECT 2.79 3.625 2.96 4.945 ;
      RECT 2.2 4.945 2.96 5.115 ;
      RECT 2.2 5.115 2.71 5.365 ;
      RECT 4.815 1.305 5.025 3.08 ;
      RECT 4.485 3.08 5.025 3.29 ;
      RECT 5.085 0.625 5.295 1.135 ;
      RECT 4.485 3.29 4.655 3.455 ;
      RECT 2.79 3.455 4.655 3.625 ;
      RECT 7.22 1.475 8.38 1.665 ;
      RECT 7.58 0.61 7.82 1.475 ;
      RECT 7.22 1.665 7.43 2.03 ;
      RECT 8.07 1.665 8.38 2.145 ;
      RECT 7.18 2.03 7.43 2.36 ;
      RECT 8.55 1.265 8.75 2.36 ;
      RECT 8.1 0.97 8.75 1.265 ;
      RECT 8.1 0.61 8.83 0.97 ;
      RECT 8.1 0.595 8.38 0.61 ;
      RECT 8.965 1.545 10.55 1.715 ;
      RECT 10.21 1.505 10.55 1.545 ;
      RECT 8.965 1.715 9.135 3.105 ;
      RECT 10.3 1.715 10.55 2.52 ;
      RECT 10.21 1.335 13.315 1.505 ;
      RECT 8.805 3.105 9.135 3.435 ;
      RECT 10.21 0.64 10.46 1.335 ;
      RECT 11.585 1.505 13.315 1.58 ;
      RECT 11.62 1.25 13.315 1.335 ;
      RECT 11.585 1.58 11.865 2.635 ;
      RECT 11.62 0.72 11.95 1.25 ;
      RECT 11.38 2.635 12.045 2.965 ;
      RECT 1.455 3.84 1.785 4.67 ;
      RECT 0.86 3.585 1.785 3.84 ;
      RECT 1.455 4.67 2.03 4.84 ;
      RECT 1.86 4.84 2.03 5.625 ;
      RECT 1.86 5.625 2.11 5.955 ;
      RECT 3.59 3.925 3.92 4.17 ;
      RECT 3.14 4.17 3.92 4.59 ;
      RECT 3.14 4.59 3.42 5.285 ;
      RECT 2.88 5.285 3.42 5.455 ;
      RECT 2.88 5.455 3.05 5.625 ;
      RECT 2.8 5.625 3.05 5.955 ;
      RECT 5.925 3.35 7.405 3.43 ;
      RECT 5.925 3.095 8.37 3.35 ;
      RECT 8.09 3.35 8.37 4.685 ;
      RECT 7.6 3.085 8.37 3.095 ;
      RECT 7.6 2.03 7.895 3.085 ;
      RECT 6.57 3.985 6.9 4.695 ;
      RECT 6.465 3.705 7.005 3.985 ;
      RECT 6.04 3.795 6.295 4.155 ;
      RECT 6.04 4.155 6.35 4.605 ;
      RECT 5.72 4.605 6.35 4.775 ;
      RECT 5.72 4.775 5.89 5.475 ;
      RECT 5.38 5.475 5.89 5.69 ;
      RECT 5.38 5.69 6.06 6.065 ;
      RECT 4.5 4.865 5.55 5.035 ;
      RECT 5.38 4.435 5.55 4.865 ;
      RECT 5.38 4.265 5.665 4.435 ;
      RECT 5.495 2.895 5.665 4.265 ;
      RECT 5.495 2.225 5.825 2.895 ;
      RECT 4.5 4.135 4.835 4.865 ;
      RECT 4.5 5.035 4.67 5.58 ;
      RECT 4.3 5.58 4.67 5.955 ;
      RECT 5.005 3.985 5.21 4.695 ;
      RECT 5.005 3.965 5.325 3.985 ;
      RECT 4.09 3.795 5.325 3.965 ;
      RECT 4.09 3.965 4.33 4.705 ;
      RECT 4.78 3.745 5.325 3.795 ;
      RECT 10.55 3.755 10.88 4.94 ;
      RECT 9.36 4.94 12.05 5.11 ;
      RECT 9.36 5.11 9.61 5.24 ;
      RECT 9.36 4.91 9.61 4.94 ;
  END
END scs8ls_lpflow_srsdfxtp2_2

MACRO scs8ls_lpflow_srsdfstp2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 16.8 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.32 1.145 5.625 1.815 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.059 LAYER li1 ;
  END SCD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.935 0.37 16.225 3.015 ;
    END
    ANTENNADIFFAREA 0.5544 ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1 ;
  END Q

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.1 4.695 1.42 5.365 ;
    END
    ANTENNAGATEAREA 0.318 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.13 LAYER li1 ;
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.145 0.455 1.815 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.3 5.205 6.61 5.875 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.06 LAYER li1 ;
  END CLK

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.64 5.6 7.81 6.235 ;
        RECT 5.305 6.235 7.81 6.405 ;
        RECT 5.305 5.525 5.475 6.235 ;
        RECT 5.145 4.885 5.475 5.525 ;
        RECT 7.64 5.535 8.485 5.6 ;
        RECT 8.3 5.205 8.89 5.43 ;
        RECT 7.64 5.43 8.89 5.535 ;
    END
    ANTENNAGATEAREA 0.598 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.191 LAYER li1 ;
  END SLEEPB

  PIN SETB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met1 ;
        RECT 2.14 2.705 15.1 2.845 ;
        RECT 14.45 2.845 15.1 2.92 ;
        RECT 14.45 2.69 15.1 2.705 ;
        RECT 2.14 2.845 2.795 2.92 ;
        RECT 8.235 2.845 8.885 2.92 ;
        RECT 2.14 2.69 2.795 2.705 ;
        RECT 8.235 2.69 8.885 2.705 ;
    END
    ANTENNAGATEAREA 0.378 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 9.121 LAYER met1 ;
  END SETB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 16.8 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 16.8 6.905 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 16.8 3.575 ;
        RECT 2.975 3.075 6.145 3.085 ;
        RECT 11.85 2.985 13.33 3.085 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 3.715 16.73 3.985 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 13.04 3.285 13.21 3.455 ;
      RECT 12.645 3.075 12.815 3.245 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 6.575 12.805 6.745 ;
      RECT 12.285 3.075 12.455 3.245 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 6.575 12.325 6.745 ;
      RECT 11.915 3.03 12.085 3.2 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 6.575 11.845 6.745 ;
      RECT 11.54 3.785 11.71 3.955 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 6.575 11.365 6.745 ;
      RECT 11.18 3.785 11.35 3.955 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 6.575 10.885 6.745 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 6.155 3.785 6.325 3.955 ;
      RECT 5.265 3.785 5.435 3.955 ;
      RECT 10.235 6.575 10.405 6.745 ;
      RECT 5.915 3.105 6.085 3.275 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 6.575 9.925 6.745 ;
      RECT 9.615 3.245 9.785 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 6.575 9.445 6.745 ;
      RECT 9.255 3.18 9.425 3.35 ;
      RECT 8.895 3.18 9.065 3.35 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 6.575 8.965 6.745 ;
      RECT 8.655 2.72 8.825 2.89 ;
      RECT 8.535 3.18 8.705 3.35 ;
      RECT 8.295 2.72 8.465 2.89 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 6.575 8.485 6.745 ;
      RECT 8.255 3.765 8.425 3.935 ;
      RECT 8.175 3.18 8.345 3.35 ;
      RECT 7.895 3.765 8.065 3.935 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 6.575 8.005 6.745 ;
      RECT 7.815 3.18 7.985 3.35 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 7.455 3.18 7.625 3.35 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 6.575 7.525 6.745 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 6.575 7.045 6.745 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.555 3.105 5.725 3.275 ;
      RECT 6.395 6.575 6.565 6.745 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.195 3.105 5.365 3.275 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 4.835 3.105 5.005 3.275 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 4.475 3.105 4.645 3.275 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 4.115 3.105 4.285 3.275 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.755 3.105 3.925 3.275 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.395 3.105 3.565 3.275 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.105 3.205 3.275 ;
      RECT 3.035 6.575 3.205 6.745 ;
      RECT 2.56 2.72 2.73 2.89 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 2.2 2.72 2.37 2.89 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 16.475 6.575 16.645 6.745 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.995 6.575 16.165 6.745 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.515 6.575 15.685 6.745 ;
      RECT 15.155 3.295 15.325 3.465 ;
      RECT 14.87 2.72 15.04 2.89 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 6.575 15.205 6.745 ;
      RECT 14.795 3.295 14.965 3.465 ;
      RECT 14.51 2.72 14.68 2.89 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 6.575 14.725 6.745 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 6.575 14.245 6.745 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 6.575 13.765 6.745 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 6.575 13.285 6.745 ;
    LAYER li1 ;
      RECT 5.645 4.865 6.695 5.035 ;
      RECT 5.645 4.125 5.975 4.865 ;
      RECT 5.92 5.035 6.13 6.01 ;
      RECT 7.465 4.155 7.795 4.525 ;
      RECT 7.465 3.795 7.72 4.155 ;
      RECT 7.01 4.525 7.795 4.695 ;
      RECT 7.01 4.695 7.18 5.475 ;
      RECT 6.82 5.475 7.18 5.69 ;
      RECT 6.82 5.69 7.47 6.065 ;
      RECT 11.915 2.87 13.305 3.245 ;
      RECT 11.915 1.895 12.295 2.87 ;
      RECT 12.94 3.245 13.305 4.065 ;
      RECT 12.94 4.065 13.415 4.395 ;
      RECT 10.46 3.605 10.96 4.685 ;
      RECT 10.745 3.585 10.96 3.605 ;
      RECT 10.46 4.685 10.63 5.69 ;
      RECT 10.745 3.415 12.77 3.585 ;
      RECT 10.46 5.69 10.8 6.02 ;
      RECT 12.49 3.585 12.77 4.305 ;
      RECT 11.13 3.755 11.79 4.685 ;
      RECT 11.99 3.755 12.32 4.875 ;
      RECT 11.99 4.875 13.465 4.91 ;
      RECT 10.8 4.91 13.465 5.11 ;
      RECT 10.8 5.11 11.05 5.24 ;
      RECT 12.47 5.11 13.465 5.19 ;
      RECT 12.47 5.19 12.705 6.02 ;
      RECT 8.525 4.155 9.36 4.865 ;
      RECT 8.6 3.795 9.36 4.155 ;
      RECT 7.365 4.865 9.36 5.035 ;
      RECT 9.03 3.73 9.36 3.795 ;
      RECT 9.06 5.035 9.36 5.38 ;
      RECT 9.06 5.38 9.91 5.55 ;
      RECT 9.06 5.55 9.23 5.705 ;
      RECT 9.74 5.55 9.91 6.19 ;
      RECT 8.77 5.705 9.23 6.065 ;
      RECT 9.74 6.19 11.34 6.39 ;
      RECT 11.17 5.55 11.34 6.19 ;
      RECT 11.17 5.38 12.3 5.55 ;
      RECT 12.13 5.55 12.3 6.19 ;
      RECT 11.225 5.285 12.3 5.38 ;
      RECT 12.13 6.19 13.445 6.39 ;
      RECT 13.135 5.525 13.445 6.19 ;
      RECT 7.365 5.035 8.035 5.26 ;
      RECT 13.975 3.745 14.345 4.275 ;
      RECT 13.975 2.65 14.265 3.745 ;
      RECT 13.975 4.275 14.915 5.16 ;
      RECT 13.975 5.16 14.235 5.33 ;
      RECT 14.745 5.16 14.915 5.72 ;
      RECT 13.615 5.33 14.235 5.66 ;
      RECT 14.745 5.72 15.095 6.05 ;
      RECT 15.15 4.23 15.4 4.775 ;
      RECT 15.15 4.775 16.3 4.945 ;
      RECT 16.07 4.23 16.3 4.775 ;
      RECT 14.51 2.455 15.04 3.125 ;
      RECT 14.435 3.295 16.8 3.415 ;
      RECT 15.475 3.245 16.8 3.295 ;
      RECT 16.395 1.855 16.685 3.245 ;
      RECT 15.57 3.575 15.9 4.605 ;
      RECT 14.435 3.415 15.9 3.575 ;
      RECT 15.475 2.19 15.765 3.245 ;
      RECT 14.435 1.84 15.765 2.19 ;
      RECT 6.38 0.255 8.73 0.425 ;
      RECT 8.56 0.425 8.73 1.03 ;
      RECT 8.56 1.03 10.455 1.125 ;
      RECT 7.925 1.125 10.455 1.2 ;
      RECT 10.285 0.425 10.455 1.03 ;
      RECT 7.925 1.2 8.73 1.295 ;
      RECT 10.285 0.255 11.82 0.425 ;
      RECT 7.925 1.295 8.515 1.455 ;
      RECT 11.65 0.425 11.82 1.11 ;
      RECT 11.65 1.11 13.09 1.345 ;
      RECT 12.835 1.345 13.09 2.31 ;
      RECT 3.85 3.615 4.02 4.945 ;
      RECT 2.825 4.945 4.02 5.115 ;
      RECT 2.825 5.115 3.335 5.365 ;
      RECT 6.38 0.425 6.63 3.445 ;
      RECT 3.85 3.445 6.63 3.615 ;
      RECT 0 -0.085 16.8 0.085 ;
      RECT 16.395 0.085 16.675 1.15 ;
      RECT 5.88 0.085 6.21 0.955 ;
      RECT 9.21 0.085 10.115 0.86 ;
      RECT 11.99 0.085 15.765 0.285 ;
      RECT 11.99 0.285 12.645 0.94 ;
      RECT 14.405 0.285 15.765 1.125 ;
      RECT 0.965 0.085 1.3 1.06 ;
      RECT 2.93 0.085 3.25 1.015 ;
      RECT 4.56 0.085 4.81 0.975 ;
      RECT 0 6.575 16.8 6.745 ;
      RECT 8.01 6.265 9.57 6.575 ;
      RECT 11.51 5.72 11.96 6.575 ;
      RECT 14.28 6.22 16.285 6.575 ;
      RECT 8.01 5.77 8.6 6.265 ;
      RECT 9.4 5.72 9.57 6.265 ;
      RECT 14.28 5.83 14.575 6.22 ;
      RECT 15.955 5.72 16.285 6.22 ;
      RECT 14.405 5.33 14.575 5.83 ;
      RECT 1.1 6.28 4.11 6.575 ;
      RECT 4.73 5.68 5.06 6.575 ;
      RECT 2.05 5.625 2.315 6.28 ;
      RECT 2.915 5.625 3.245 6.28 ;
      RECT 3.845 5.625 4.11 6.28 ;
      RECT 1.1 5.605 1.395 6.28 ;
      RECT 4.98 0.645 5.6 0.975 ;
      RECT 3.975 1.32 4.225 1.815 ;
      RECT 3.975 1.145 5.15 1.32 ;
      RECT 4.85 1.32 5.1 2.655 ;
      RECT 4.98 0.975 5.15 1.145 ;
      RECT 3.585 0.975 3.805 1.985 ;
      RECT 3.45 0.255 4.1 0.975 ;
      RECT 3.585 1.985 4.14 2.205 ;
      RECT 3.91 2.205 4.14 2.655 ;
      RECT 2.495 1.185 3.415 1.855 ;
      RECT 2.495 0.65 2.76 1.185 ;
      RECT 2.495 1.855 2.76 2.34 ;
      RECT 1.97 0.975 2.19 1.99 ;
      RECT 1.675 0.255 2.325 0.975 ;
      RECT 1.515 1.99 2.19 2.175 ;
      RECT 1.515 2.175 1.785 2.66 ;
      RECT 0.625 1.615 1.8 1.82 ;
      RECT 1.55 1.145 1.8 1.615 ;
      RECT 0.625 0.975 0.795 1.615 ;
      RECT 0.625 1.82 0.845 2.66 ;
      RECT 0.095 0.645 0.795 0.975 ;
      RECT 7.575 1.71 9.615 1.88 ;
      RECT 7.575 1.185 7.755 1.71 ;
      RECT 8.28 1.88 8.49 2.345 ;
      RECT 9.345 1.88 9.615 2.335 ;
      RECT 7.305 0.955 7.755 1.185 ;
      RECT 7.305 0.595 8.39 0.955 ;
      RECT 10.585 1.59 10.895 2.38 ;
      RECT 10.045 1.54 10.895 1.59 ;
      RECT 9.065 1.37 10.895 1.54 ;
      RECT 10.625 0.625 10.895 1.37 ;
      RECT 11.145 1.515 12.665 1.725 ;
      RECT 11.145 0.595 11.48 1.515 ;
      RECT 11.145 1.725 11.46 3.025 ;
      RECT 12.465 1.725 12.665 2.48 ;
      RECT 10.225 3.025 11.46 3.245 ;
      RECT 12.465 2.48 13.805 2.7 ;
      RECT 10.225 3.245 10.575 3.435 ;
      RECT 13.26 1.625 13.805 2.48 ;
      RECT 13.475 2.7 13.805 3.68 ;
      RECT 13.26 1.295 15.765 1.625 ;
      RECT 13.26 0.755 13.97 1.295 ;
      RECT 0 3.245 1.345 3.415 ;
      RECT 0.095 2.84 1.345 3.245 ;
      RECT 1.015 1.99 1.345 2.84 ;
      RECT 0.16 3.415 0.52 4.84 ;
      RECT 0.095 2.02 0.455 2.84 ;
      RECT 2.895 3.275 3.265 4.775 ;
      RECT 2.895 3.24 6.21 3.275 ;
      RECT 2.93 2.855 6.21 3.24 ;
      RECT 2.93 2.025 3.28 2.855 ;
      RECT 4.315 2.835 6.21 2.855 ;
      RECT 5.27 2.015 6.21 2.835 ;
      RECT 4.315 1.985 4.68 2.835 ;
      RECT 4.215 3.925 4.995 4.595 ;
      RECT 4.215 4.595 4.54 5.285 ;
      RECT 3.505 5.285 4.54 5.455 ;
      RECT 3.505 5.455 3.675 5.535 ;
      RECT 4.28 5.455 4.54 5.955 ;
      RECT 3.415 5.535 3.675 5.955 ;
      RECT 2.14 2.61 2.76 2.94 ;
      RECT 1.59 3.84 1.99 4.64 ;
      RECT 0.895 3.585 1.99 3.84 ;
      RECT 1.59 4.64 2.655 4.84 ;
      RECT 1.59 4.84 1.88 5.955 ;
      RECT 2.485 4.84 2.655 5.535 ;
      RECT 2.485 5.535 2.745 5.955 ;
      RECT 0.69 4.17 0.93 5.255 ;
      RECT 0.235 5.255 0.93 5.955 ;
      RECT 7.365 3.09 9.81 3.535 ;
      RECT 9.53 3.535 9.81 4.685 ;
      RECT 9.005 2.855 9.81 3.09 ;
      RECT 9.005 2.505 10.385 2.855 ;
      RECT 9.005 2.345 9.175 2.505 ;
      RECT 10.045 1.99 10.385 2.505 ;
      RECT 8.66 2.05 9.175 2.345 ;
      RECT 8.245 2.54 8.835 2.92 ;
      RECT 7.965 3.985 8.355 4.695 ;
      RECT 7.89 3.705 8.43 3.985 ;
      RECT 5.235 3.955 5.475 4.715 ;
      RECT 5.235 3.785 6.355 3.955 ;
      RECT 6.145 3.955 6.355 4.695 ;
      RECT 6.525 4.23 6.695 4.865 ;
      RECT 6.525 4.06 6.97 4.23 ;
      RECT 6.8 2.895 6.97 4.06 ;
      RECT 6.8 2.225 7.13 2.895 ;
  END
END scs8ls_lpflow_srsdfstp2_2

MACRO scs8ls_lpflow_srsdfrtp2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 17.28 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.5 1.125 6.085 1.44 ;
        RECT 5.5 1.44 5.725 1.795 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.183 LAYER li1 ;
  END SCD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.415 0.37 16.705 3.015 ;
    END
    ANTENNADIFFAREA 0.5544 ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1 ;
  END Q

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.49 5.035 2.08 5.455 ;
    END
    ANTENNAGATEAREA 0.318 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.134 LAYER li1 ;
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.095 0.425 1.765 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.058 LAYER li1 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.68 4.895 7.195 5.515 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.091 LAYER li1 ;
  END CLK

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.15 5.205 9.85 5.38 ;
        RECT 8.615 5.38 9.85 5.535 ;
        RECT 8.615 5.535 9.32 5.55 ;
        RECT 8.615 5.55 8.785 6.235 ;
        RECT 7.225 6.235 8.785 6.405 ;
        RECT 7.225 6.205 7.595 6.235 ;
        RECT 7.425 5.265 7.595 6.205 ;
        RECT 7.425 4.935 7.74 5.265 ;
    END
    ANTENNAGATEAREA 0.598 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.986 LAYER li1 ;
  END SLEEPB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 17.28 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 17.28 6.905 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 17.28 3.575 ;
        RECT 6.38 2.985 8.11 3.085 ;
        RECT 10.405 2.985 15.03 3.085 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 3.715 17.21 3.985 ;
    END
  END kapwr

  PIN RESETB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met1 ;
        RECT 2.535 2.705 15.83 2.845 ;
        RECT 15.17 2.845 15.83 2.935 ;
        RECT 15.515 2.69 15.83 2.705 ;
        RECT 2.535 2.845 3.215 2.935 ;
        RECT 8.45 2.845 9.1 2.92 ;
        RECT 2.535 2.69 3.215 2.705 ;
        RECT 8.45 2.69 9.1 2.705 ;
    END
    ANTENNAGATEAREA 0.378 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 9.3765 LAYER met1 ;
  END RESETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 8.87 2.72 9.04 2.89 ;
      RECT 8.855 3.765 9.025 3.935 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 6.575 8.965 6.745 ;
      RECT 8.51 2.72 8.68 2.89 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 6.575 8.485 6.745 ;
      RECT 8.04 3.785 8.21 3.955 ;
      RECT 7.88 3.105 8.05 3.275 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 6.575 8.005 6.745 ;
      RECT 7.68 3.785 7.85 3.955 ;
      RECT 7.52 3.105 7.69 3.275 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 6.575 7.525 6.745 ;
      RECT 7.16 3.105 7.33 3.275 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 6.575 7.045 6.745 ;
      RECT 6.8 3.105 6.97 3.275 ;
      RECT 6.795 3.785 6.965 3.955 ;
      RECT 6.44 3.015 6.61 3.185 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 6.575 6.565 6.745 ;
      RECT 6.315 3.375 6.485 3.545 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 5.475 3.245 5.645 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 5.105 3.245 5.275 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 4.525 3.245 4.695 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 4.155 3.245 4.325 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 3.785 3.245 3.955 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 3.415 3.245 3.585 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 6.575 3.205 6.745 ;
      RECT 2.985 2.735 3.155 2.905 ;
      RECT 2.595 2.735 2.765 2.905 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 16.995 3.245 17.165 3.415 ;
      RECT 16.955 -0.085 17.125 0.085 ;
      RECT 16.955 6.575 17.125 6.745 ;
      RECT 16.635 3.245 16.805 3.415 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 16.475 6.575 16.645 6.745 ;
      RECT 16.275 3.295 16.445 3.465 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 6.575 16.165 6.745 ;
      RECT 15.915 3.295 16.085 3.465 ;
      RECT 15.6 2.735 15.77 2.905 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 6.575 15.685 6.745 ;
      RECT 15.24 2.735 15.41 2.905 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 6.575 15.205 6.745 ;
      RECT 14.8 3.015 14.97 3.185 ;
      RECT 14.8 3.375 14.97 3.545 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 6.575 14.725 6.745 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 6.575 14.245 6.745 ;
      RECT 13.95 3.015 14.12 3.185 ;
      RECT 13.95 3.375 14.12 3.545 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 6.575 13.765 6.745 ;
      RECT 13.59 3.015 13.76 3.185 ;
      RECT 13.23 3.015 13.4 3.185 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 6.575 13.285 6.745 ;
      RECT 12.87 3.015 13.04 3.185 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 1.26 3.245 1.43 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 0.89 3.245 1.06 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 0.525 3.245 0.695 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 6.575 12.805 6.745 ;
      RECT 12.51 3.015 12.68 3.185 ;
      RECT 12.5 3.785 12.67 3.955 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 6.575 12.325 6.745 ;
      RECT 12.14 3.785 12.31 3.955 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 6.575 11.845 6.745 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 6.575 11.365 6.745 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 6.575 10.885 6.745 ;
      RECT 10.51 3.375 10.68 3.545 ;
      RECT 10.465 3.015 10.635 3.185 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 6.575 10.405 6.745 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 6.575 9.925 6.745 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 6.575 9.445 6.745 ;
      RECT 9.215 3.765 9.385 3.935 ;
    LAYER li1 ;
      RECT 9.485 4.155 9.815 4.865 ;
      RECT 9.99 3.52 10.32 3.795 ;
      RECT 8.81 4.865 10.19 4.955 ;
      RECT 8.31 4.955 10.19 5.035 ;
      RECT 10.02 5.035 10.19 5.38 ;
      RECT 10.02 5.38 11.22 5.55 ;
      RECT 10.02 5.55 10.19 5.735 ;
      RECT 11.05 5.55 11.22 6.22 ;
      RECT 9.825 5.735 10.19 6.065 ;
      RECT 11.05 6.22 12.3 6.39 ;
      RECT 12.13 5.55 12.3 6.22 ;
      RECT 12.13 5.38 13.26 5.55 ;
      RECT 13.09 5.55 13.26 6.22 ;
      RECT 12.345 5.285 12.675 5.38 ;
      RECT 13.09 6.22 14.425 6.39 ;
      RECT 14.095 5.865 14.425 6.22 ;
      RECT 14.095 5.525 14.405 5.865 ;
      RECT 8.31 5.035 8.98 5.21 ;
      RECT 8.51 3.135 10.15 3.305 ;
      RECT 9.98 1.8 10.15 3.135 ;
      RECT 9.98 1.63 11.22 1.8 ;
      RECT 10.94 1.8 11.22 2.69 ;
      RECT 6.34 5.685 7.255 6.015 ;
      RECT 6.18 4.725 6.51 5.21 ;
      RECT 6.34 5.21 6.51 5.685 ;
      RECT 7.215 3.705 7.465 4.555 ;
      RECT 7.295 3.615 7.465 3.705 ;
      RECT 6.18 4.555 7.465 4.725 ;
      RECT 7.295 3.445 8.68 3.615 ;
      RECT 8.51 3.305 8.68 3.445 ;
      RECT 8.955 3.985 9.285 4.695 ;
      RECT 8.85 3.705 9.39 3.985 ;
      RECT 8.41 2.655 9.14 2.93 ;
      RECT 8.41 1.935 9.08 2.655 ;
      RECT 8.425 3.795 8.68 4.155 ;
      RECT 8.425 4.155 8.755 4.615 ;
      RECT 7.97 4.615 8.755 4.695 ;
      RECT 7.97 4.695 8.595 4.785 ;
      RECT 7.97 4.785 8.14 5.475 ;
      RECT 7.765 5.475 8.14 5.735 ;
      RECT 7.765 5.735 8.445 6.065 ;
      RECT 7.635 3.785 8.255 4.445 ;
      RECT 6.275 3.275 6.525 4.385 ;
      RECT 6.275 3.085 8.15 3.275 ;
      RECT 6.275 1.95 6.69 3.085 ;
      RECT 7.855 1.93 8.15 3.085 ;
      RECT 6.715 3.705 7.045 4.385 ;
      RECT 12.95 3.755 13.28 4.94 ;
      RECT 11.76 4.94 14.855 5.11 ;
      RECT 11.76 5.11 12.01 5.24 ;
      RECT 13.45 5.11 13.7 6.05 ;
      RECT 11.76 4.91 12.01 4.94 ;
      RECT 14.265 5.11 14.855 5.16 ;
      RECT 14.265 4.83 14.855 4.94 ;
      RECT 12.45 2.955 14.17 3.245 ;
      RECT 12.45 1.945 13.03 2.955 ;
      RECT 13.9 3.245 14.17 4.165 ;
      RECT 12.745 1.825 13.03 1.945 ;
      RECT 13.9 4.165 14.455 4.445 ;
      RECT 11.42 3.585 11.795 4.685 ;
      RECT 11.42 3.415 13.73 3.585 ;
      RECT 11.42 4.685 11.59 5.72 ;
      RECT 13.45 3.585 13.73 4.305 ;
      RECT 11.42 5.72 11.76 6.05 ;
      RECT 12.42 3.985 12.75 4.685 ;
      RECT 12.09 3.755 12.75 3.985 ;
      RECT 10.49 3.4 10.78 4.685 ;
      RECT 10.49 3.35 10.695 3.4 ;
      RECT 10.405 2.73 10.695 3.35 ;
      RECT 10.405 1.97 10.77 2.73 ;
      RECT 15.18 2.935 15.43 3.4 ;
      RECT 15.18 2.705 15.83 2.935 ;
      RECT 15.025 4.995 16.955 5.165 ;
      RECT 16.625 5.165 16.955 6.05 ;
      RECT 16.45 4.275 16.78 4.995 ;
      RECT 14.66 4.045 15.265 4.215 ;
      RECT 14.66 3.995 14.91 4.045 ;
      RECT 15.025 4.215 15.265 4.995 ;
      RECT 14.34 3.745 14.91 3.995 ;
      RECT 14.34 2.88 14.59 3.745 ;
      RECT 15.025 5.165 15.195 5.33 ;
      RECT 14.575 5.33 15.195 5.5 ;
      RECT 14.575 5.5 14.825 5.685 ;
      RECT 14.76 2.25 15.01 3.575 ;
      RECT 14.505 1.92 15.01 2.25 ;
      RECT 15.6 3.415 16.75 4.075 ;
      RECT 15.6 3.245 17.28 3.415 ;
      RECT 15.6 3.185 17.145 3.245 ;
      RECT 16.875 1.855 17.145 3.185 ;
      RECT 15.6 4.075 15.93 4.605 ;
      RECT 16 1.855 16.245 3.185 ;
      RECT 1.08 5.925 1.32 5.955 ;
      RECT 0.6 5.255 1.32 5.925 ;
      RECT 1.08 4.17 1.32 5.255 ;
      RECT 0 6.575 17.28 6.745 ;
      RECT 8.955 5.72 9.285 6.575 ;
      RECT 10.36 5.72 10.75 6.575 ;
      RECT 12.5 5.72 12.89 6.575 ;
      RECT 15.365 5.72 16.085 6.575 ;
      RECT 15.365 5.355 15.615 5.72 ;
      RECT 1.51 5.625 1.775 6.575 ;
      RECT 2.64 5.77 2.97 6.575 ;
      RECT 4.37 5.77 4.7 6.575 ;
      RECT 5.84 5.67 6.17 6.575 ;
      RECT 3.505 5.625 3.835 6.575 ;
      RECT 0 -0.085 17.28 0.085 ;
      RECT 16.875 0.085 17.175 1.15 ;
      RECT 6.02 0.085 6.35 0.86 ;
      RECT 8.115 0.085 8.325 0.94 ;
      RECT 10.415 0.085 11.825 0.97 ;
      RECT 14.945 0.085 15.195 0.81 ;
      RECT 15.965 0.085 16.245 1.15 ;
      RECT 1.03 0.085 1.36 0.97 ;
      RECT 3.085 0.085 3.405 0.99 ;
      RECT 4.615 0.085 4.935 1 ;
      RECT 1.74 0.57 2.39 0.895 ;
      RECT 2.115 0.895 2.39 0.925 ;
      RECT 2.14 0.255 2.39 0.57 ;
      RECT 2.115 0.925 2.325 1.935 ;
      RECT 1.62 1.935 2.325 2.145 ;
      RECT 1.62 2.145 1.91 2.605 ;
      RECT 0.69 1.35 0.91 2.605 ;
      RECT 0.69 1.18 1.945 1.35 ;
      RECT 1.615 1.35 1.945 1.735 ;
      RECT 1.615 1.125 1.945 1.18 ;
      RECT 0.69 0.925 0.86 1.18 ;
      RECT 0.16 0.595 0.86 0.925 ;
      RECT 2.495 1.095 2.915 1.825 ;
      RECT 2.645 0.64 2.915 1.095 ;
      RECT 2.66 1.825 2.915 2.34 ;
      RECT 5.105 0.625 5.805 0.955 ;
      RECT 4.02 1.415 5.33 1.63 ;
      RECT 4.02 1.125 4.35 1.415 ;
      RECT 5.105 0.955 5.33 1.415 ;
      RECT 4.02 1.63 4.35 1.735 ;
      RECT 4.975 1.63 5.215 2.605 ;
      RECT 3.64 0.925 3.85 1.935 ;
      RECT 3.575 0.6 4.225 0.925 ;
      RECT 3.64 1.935 4.265 2.145 ;
      RECT 3.575 0.255 3.825 0.6 ;
      RECT 4.055 2.145 4.265 2.605 ;
      RECT 8.495 0.255 10.245 0.425 ;
      RECT 10.075 0.425 10.245 1.15 ;
      RECT 10.075 1.15 12.165 1.32 ;
      RECT 10.075 1.32 10.925 1.46 ;
      RECT 11.995 0.425 12.165 1.15 ;
      RECT 11.995 0.255 13.445 0.425 ;
      RECT 13.275 0.425 13.445 0.465 ;
      RECT 13.275 0.465 13.555 1.135 ;
      RECT 6.52 0.425 6.69 1.61 ;
      RECT 5.895 1.61 6.69 1.78 ;
      RECT 5.895 1.78 6.105 3.585 ;
      RECT 4.035 3.585 6.105 3.755 ;
      RECT 5.775 3.755 6.105 4.155 ;
      RECT 5.71 4.155 6.105 4.365 ;
      RECT 5.71 4.365 5.92 5.29 ;
      RECT 5.46 5.29 5.92 5.5 ;
      RECT 5.46 5.5 5.67 6.02 ;
      RECT 4.035 3.755 4.205 4.945 ;
      RECT 3.335 4.945 4.205 5.115 ;
      RECT 3.335 5.115 4.005 5.26 ;
      RECT 7.775 0.425 7.945 1.12 ;
      RECT 6.52 0.255 7.945 0.425 ;
      RECT 7.775 1.12 8.665 1.29 ;
      RECT 8.495 0.425 8.665 1.12 ;
      RECT 9.38 1.305 9.55 1.93 ;
      RECT 9.19 0.94 9.55 1.305 ;
      RECT 9.25 1.93 9.55 2.26 ;
      RECT 8.835 0.595 9.905 0.94 ;
      RECT 7.395 1.475 9.21 1.665 ;
      RECT 7.395 0.61 7.605 1.475 ;
      RECT 7.395 1.665 7.655 2.26 ;
      RECT 8.54 1.665 9.21 1.725 ;
      RECT 6.86 0.61 7.1 2.645 ;
      RECT 6.86 2.645 7.685 2.895 ;
      RECT 11.85 1.49 12.575 1.775 ;
      RECT 12.335 1.475 12.575 1.49 ;
      RECT 11.85 1.775 12.18 2.9 ;
      RECT 12.335 1.305 13.975 1.475 ;
      RECT 10.865 2.9 12.18 3.07 ;
      RECT 12.335 0.625 12.575 1.305 ;
      RECT 13.675 1.475 13.975 1.56 ;
      RECT 13.725 0.48 13.975 1.305 ;
      RECT 10.865 3.07 11.455 3.23 ;
      RECT 13.675 1.56 16.245 1.65 ;
      RECT 15.655 1.32 16.245 1.56 ;
      RECT 13.675 1.65 15.825 1.73 ;
      RECT 13.675 1.73 13.965 2.295 ;
      RECT 15.375 1.73 15.665 2.295 ;
      RECT 14.475 0.98 15.625 1.15 ;
      RECT 14.475 0.48 14.775 0.98 ;
      RECT 15.365 0.48 15.625 0.98 ;
      RECT 0.505 4.11 0.87 4.84 ;
      RECT 0.505 3.415 0.725 4.11 ;
      RECT 0 3.245 1.46 3.415 ;
      RECT 0.22 2.79 1.46 3.245 ;
      RECT 0.22 2.785 1.41 2.79 ;
      RECT 0.22 1.935 0.5 2.785 ;
      RECT 1.08 1.935 1.41 2.785 ;
      RECT 0.925 3.585 2.61 3.84 ;
      RECT 2.25 3.84 2.61 4.845 ;
      RECT 2.25 4.845 2.46 5.43 ;
      RECT 2.25 5.43 3.335 5.6 ;
      RECT 2.25 5.6 2.46 5.955 ;
      RECT 3.145 5.6 3.335 5.995 ;
      RECT 3.505 3.415 3.835 4.775 ;
      RECT 3.355 2.79 5.725 3.415 ;
      RECT 3.355 2.525 3.825 2.79 ;
      RECT 5.385 1.97 5.725 2.79 ;
      RECT 4.475 1.935 4.805 2.79 ;
      RECT 3.115 2.315 3.825 2.525 ;
      RECT 3.115 1.925 3.445 2.315 ;
      RECT 5.21 3.925 5.54 4.17 ;
      RECT 4.77 4.17 5.54 4.595 ;
      RECT 4.77 4.595 5.09 5.43 ;
      RECT 4.005 5.43 5.13 5.6 ;
      RECT 4.005 5.6 4.195 5.995 ;
      RECT 4.88 5.6 5.13 5.955 ;
      RECT 2.565 2.695 3.185 3.025 ;
      RECT 9.56 4.11 9.815 4.155 ;
      RECT 9.56 3.795 10.32 4.11 ;
  END
END scs8ls_lpflow_srsdfrtp2_2

MACRO scs8ls_lpflow_srsdfxtp2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 14.88 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.47 4.305 1.795 ;
        RECT 4.025 1.125 4.305 1.47 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.134 LAYER li1 ;
  END SCD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.555 0.37 13.845 3.015 ;
    END
    ANTENNADIFFAREA 0.5097 ;
    ANTENNAPARTIALMETALSIDEAREA 0.519 LAYER li1 ;
  END Q

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045 5.035 1.69 5.455 ;
    END
    ANTENNAGATEAREA 0.318 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.145 LAYER li1 ;
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.095 0.455 1.765 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.84 5.205 5.17 5.875 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END CLK

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.86 5.205 7.45 5.445 ;
        RECT 6.23 5.445 7.45 5.535 ;
        RECT 6.23 5.535 7.015 5.615 ;
        RECT 6.23 5.615 6.4 6.235 ;
        RECT 3.72 6.235 6.4 6.405 ;
        RECT 3.72 5.455 3.95 6.235 ;
        RECT 3.59 5.225 3.95 5.455 ;
        RECT 3.59 4.8 3.92 5.225 ;
    END
    ANTENNAGATEAREA 0.598 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.231 LAYER li1 ;
  END SLEEPB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.88 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 14.88 6.905 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.88 3.575 ;
        RECT 9.295 2.985 9.945 3.085 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 3.715 14.81 3.985 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 6.575 9.445 6.745 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 6.575 8.965 6.745 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 6.575 8.485 6.745 ;
      RECT 8.175 3.245 8.345 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 6.575 8.005 6.745 ;
      RECT 7.815 3.18 7.985 3.35 ;
      RECT 7.455 3.18 7.625 3.35 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 6.575 14.725 6.745 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 6.575 7.525 6.745 ;
      RECT 7.095 3.18 7.265 3.35 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 6.575 7.045 6.745 ;
      RECT 6.825 3.765 6.995 3.935 ;
      RECT 6.735 3.18 6.905 3.35 ;
      RECT 6.465 3.765 6.635 3.935 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 6.575 6.565 6.745 ;
      RECT 6.375 3.18 6.545 3.35 ;
      RECT 6.015 3.18 6.185 3.35 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 13.115 6.575 13.285 6.745 ;
      RECT 5.155 3.745 5.325 3.915 ;
      RECT 12.795 3.27 12.965 3.44 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 4.795 3.785 4.965 3.955 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 4.115 3.115 4.285 3.285 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 3.755 3.115 3.925 3.285 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 13.875 3.27 14.045 3.44 ;
      RECT 3.395 3.115 3.565 3.285 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 13.515 3.27 13.685 3.44 ;
      RECT 3.035 3.115 3.205 3.285 ;
      RECT 3.035 6.575 3.205 6.745 ;
      RECT 13.595 6.575 13.765 6.745 ;
      RECT 2.675 3.115 2.845 3.285 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 13.155 3.27 13.325 3.44 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 2.315 3.115 2.485 3.285 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 14.075 6.575 14.245 6.745 ;
      RECT 1.955 3.245 2.125 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 6.575 12.805 6.745 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 6.575 12.325 6.745 ;
      RECT 11.9 3.345 12.07 3.515 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 6.575 11.845 6.745 ;
      RECT 11.54 3.345 11.71 3.515 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 6.575 11.365 6.745 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 6.575 10.885 6.745 ;
      RECT 14.235 3.27 14.405 3.44 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 6.575 10.405 6.745 ;
      RECT 14.595 3.245 14.765 3.415 ;
      RECT 10.1 3.785 10.27 3.955 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 9.755 6.575 9.925 6.745 ;
      RECT 9.74 3.785 9.91 3.955 ;
      RECT 9.715 3.03 9.885 3.2 ;
      RECT 9.355 3.03 9.525 3.2 ;
    LAYER li1 ;
      RECT 9.36 4.91 9.61 4.94 ;
      RECT 11.05 5.11 11.3 6.02 ;
      RECT 11.72 5.11 12.05 5.19 ;
      RECT 11.72 4.875 12.05 4.94 ;
      RECT 9.02 3.775 9.395 4.685 ;
      RECT 9.02 3.605 9.475 3.775 ;
      RECT 9.02 4.685 9.19 5.69 ;
      RECT 9.305 3.585 9.475 3.605 ;
      RECT 9.02 5.69 9.36 6.02 ;
      RECT 9.305 3.415 11.22 3.585 ;
      RECT 11.05 3.585 11.22 3.635 ;
      RECT 11.05 3.635 11.33 4.305 ;
      RECT 9.305 2.985 9.935 3.245 ;
      RECT 9.41 1.885 9.74 2.985 ;
      RECT 7.1 4.155 7.43 4.865 ;
      RECT 7.175 4.11 7.43 4.155 ;
      RECT 6.52 4.865 7.79 4.945 ;
      RECT 7.175 3.795 7.92 4.11 ;
      RECT 6.06 4.945 7.79 5.035 ;
      RECT 7.575 3.52 7.92 3.795 ;
      RECT 7.62 5.035 7.79 5.35 ;
      RECT 7.62 5.35 8.47 5.52 ;
      RECT 7.62 5.52 7.79 5.705 ;
      RECT 8.3 5.52 8.47 6.19 ;
      RECT 7.44 5.705 7.79 6.035 ;
      RECT 8.3 6.19 9.9 6.39 ;
      RECT 9.73 5.55 9.9 6.19 ;
      RECT 9.73 5.38 10.87 5.55 ;
      RECT 10.7 5.55 10.87 6.19 ;
      RECT 9.945 5.285 10.275 5.38 ;
      RECT 10.7 6.19 12.025 6.39 ;
      RECT 11.695 5.865 12.025 6.19 ;
      RECT 11.695 5.525 12.005 5.865 ;
      RECT 6.06 5.035 6.69 5.275 ;
      RECT 10.02 3.985 10.35 4.685 ;
      RECT 9.69 3.755 10.35 3.985 ;
      RECT 12.76 3.415 14.5 3.465 ;
      RECT 12.76 3.245 14.88 3.415 ;
      RECT 13.2 3.5 13.53 4.605 ;
      RECT 12.76 3.465 13.53 3.5 ;
      RECT 12.76 2.25 13.345 3.245 ;
      RECT 12.415 1.92 13.345 2.25 ;
      RECT 13.095 1.855 13.345 1.92 ;
      RECT 11.725 3.57 12.11 4.4 ;
      RECT 11.5 3.305 12.11 3.57 ;
      RECT 12.585 4.985 14.555 5.155 ;
      RECT 14.225 5.155 14.555 6.05 ;
      RECT 14.05 4.275 14.38 4.985 ;
      RECT 12.585 3.87 12.825 4.985 ;
      RECT 12.28 3.67 12.825 3.87 ;
      RECT 12.28 2.635 12.59 3.67 ;
      RECT 12.585 5.155 12.755 5.33 ;
      RECT 12.175 5.33 12.755 5.5 ;
      RECT 12.175 5.5 12.425 5.685 ;
      RECT 0 -0.085 14.88 0.085 ;
      RECT 0.965 0.085 1.215 1.01 ;
      RECT 3.265 0.085 3.515 0.96 ;
      RECT 4.585 0.085 4.915 0.955 ;
      RECT 6.74 0.085 7.07 0.965 ;
      RECT 9.34 0.085 9.66 0.97 ;
      RECT 12.38 0.085 13.385 1.07 ;
      RECT 0 3.245 4.315 3.285 ;
      RECT 1.015 3.085 4.315 3.245 ;
      RECT 3.055 2.775 4.315 3.085 ;
      RECT 3.975 2.615 4.315 2.775 ;
      RECT 3.975 1.965 4.645 2.615 ;
      RECT 0 3.285 2.62 3.415 ;
      RECT 0.095 1.935 0.425 3.245 ;
      RECT 0.095 3.415 0.425 4.84 ;
      RECT 2.29 3.415 2.62 4.775 ;
      RECT 1.015 1.905 1.345 3.085 ;
      RECT 3.055 1.935 3.385 2.775 ;
      RECT 0 6.575 14.88 6.745 ;
      RECT 6.57 5.785 6.9 6.575 ;
      RECT 10.16 5.72 10.53 6.575 ;
      RECT 7.96 5.69 8.13 6.575 ;
      RECT 12.925 5.72 13.685 6.575 ;
      RECT 12.925 5.355 13.215 5.72 ;
      RECT 1.065 5.625 1.68 6.575 ;
      RECT 2.29 5.625 2.62 6.575 ;
      RECT 3.22 5.625 3.55 6.575 ;
      RECT 3.685 0.625 4.305 0.955 ;
      RECT 2.6 1.3 2.93 1.765 ;
      RECT 2.6 1.13 3.855 1.3 ;
      RECT 2.6 1.125 2.93 1.13 ;
      RECT 3.555 1.3 3.795 2.605 ;
      RECT 3.685 0.955 3.855 1.13 ;
      RECT 2.135 0.925 2.345 1.905 ;
      RECT 1.675 0.6 2.805 0.925 ;
      RECT 1.555 1.905 2.345 1.935 ;
      RECT 2.075 0.255 2.405 0.6 ;
      RECT 1.555 1.935 2.845 2.18 ;
      RECT 1.555 2.18 1.765 2.575 ;
      RECT 2.635 2.18 2.845 2.605 ;
      RECT 0.625 1.35 0.845 2.575 ;
      RECT 0.625 1.18 1.88 1.35 ;
      RECT 1.55 1.35 1.88 1.735 ;
      RECT 1.55 1.095 1.88 1.18 ;
      RECT 0.625 0.925 0.795 1.18 ;
      RECT 0.095 0.595 0.795 0.925 ;
      RECT 4.815 1.135 7.41 1.305 ;
      RECT 7.24 0.425 7.41 1.135 ;
      RECT 7.24 0.255 9.17 0.425 ;
      RECT 9 0.425 9.17 1.14 ;
      RECT 9 1.14 10 1.31 ;
      RECT 9.165 1.31 9.835 1.375 ;
      RECT 9.83 0.425 10 1.14 ;
      RECT 9.83 0.255 11.155 0.425 ;
      RECT 10.985 0.425 11.155 0.465 ;
      RECT 10.985 0.465 11.295 1.135 ;
      RECT 2.79 3.625 2.96 4.945 ;
      RECT 2.2 4.945 2.96 5.115 ;
      RECT 2.2 5.115 2.71 5.365 ;
      RECT 4.815 1.305 5.025 3.08 ;
      RECT 4.485 3.08 5.025 3.29 ;
      RECT 5.085 0.625 5.295 1.135 ;
      RECT 4.485 3.29 4.655 3.455 ;
      RECT 2.79 3.455 4.655 3.625 ;
      RECT 7.22 1.475 8.38 1.665 ;
      RECT 7.58 0.61 7.82 1.475 ;
      RECT 7.22 1.665 7.43 2.03 ;
      RECT 8.07 1.665 8.38 2.145 ;
      RECT 7.18 2.03 7.43 2.36 ;
      RECT 8.55 1.265 8.75 2.36 ;
      RECT 8.1 0.97 8.75 1.265 ;
      RECT 8.1 0.61 8.83 0.97 ;
      RECT 8.1 0.595 8.38 0.61 ;
      RECT 8.965 1.545 10.55 1.715 ;
      RECT 10.21 1.505 10.55 1.545 ;
      RECT 8.965 1.715 9.135 3.105 ;
      RECT 10.3 1.715 10.55 2.52 ;
      RECT 10.21 1.335 13.315 1.505 ;
      RECT 8.805 3.105 9.135 3.435 ;
      RECT 10.21 0.64 10.46 1.335 ;
      RECT 11.585 1.505 13.315 1.58 ;
      RECT 11.62 1.25 13.315 1.335 ;
      RECT 11.585 1.58 11.865 2.635 ;
      RECT 11.62 0.72 11.95 1.25 ;
      RECT 11.38 2.635 12.045 2.965 ;
      RECT 1.455 3.84 1.785 4.67 ;
      RECT 0.86 3.585 1.785 3.84 ;
      RECT 1.455 4.67 2.03 4.84 ;
      RECT 1.86 4.84 2.03 5.625 ;
      RECT 1.86 5.625 2.11 5.955 ;
      RECT 0.595 4.17 0.805 5.255 ;
      RECT 0.155 5.255 0.805 5.955 ;
      RECT 3.14 4.17 3.92 4.59 ;
      RECT 3.59 3.925 3.92 4.17 ;
      RECT 3.14 4.59 3.42 5.285 ;
      RECT 2.88 5.285 3.42 5.455 ;
      RECT 2.88 5.455 3.05 5.625 ;
      RECT 2.8 5.625 3.05 5.955 ;
      RECT 5.925 3.35 7.405 3.43 ;
      RECT 5.925 3.095 8.37 3.35 ;
      RECT 8.09 3.35 8.37 4.685 ;
      RECT 7.6 3.085 8.37 3.095 ;
      RECT 7.6 2.03 7.895 3.085 ;
      RECT 6.57 3.985 6.9 4.695 ;
      RECT 6.465 3.705 7.005 3.985 ;
      RECT 6.04 4.155 6.35 4.605 ;
      RECT 6.04 3.795 6.295 4.155 ;
      RECT 5.72 4.605 6.35 4.775 ;
      RECT 5.72 4.775 5.89 5.475 ;
      RECT 5.38 5.475 5.89 5.69 ;
      RECT 5.38 5.69 6.06 6.065 ;
      RECT 4.5 4.865 5.55 5.035 ;
      RECT 5.38 4.435 5.55 4.865 ;
      RECT 5.38 4.265 5.665 4.435 ;
      RECT 5.495 2.895 5.665 4.265 ;
      RECT 5.495 2.225 5.825 2.895 ;
      RECT 4.5 4.135 4.835 4.865 ;
      RECT 4.5 5.035 4.67 5.58 ;
      RECT 4.3 5.58 4.67 5.955 ;
      RECT 5.005 3.985 5.21 4.695 ;
      RECT 5.005 3.965 5.325 3.985 ;
      RECT 4.09 3.795 5.325 3.965 ;
      RECT 4.09 3.965 4.33 4.705 ;
      RECT 4.78 3.745 5.325 3.795 ;
      RECT 10.55 3.755 10.88 4.94 ;
      RECT 9.36 4.94 12.05 5.11 ;
      RECT 9.36 5.11 9.61 5.24 ;
  END
END scs8ls_lpflow_srsdfxtp2_1

MACRO scs8ls_lpflow_srsdfstp2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 16.8 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.32 1.145 5.625 1.815 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.059 LAYER li1 ;
  END SCD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.995 0.37 16.29 3.015 ;
    END
    ANTENNADIFFAREA 0.5097 ;
    ANTENNAPARTIALMETALSIDEAREA 0.52 LAYER li1 ;
  END Q

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.1 4.695 1.42 5.365 ;
    END
    ANTENNAGATEAREA 0.318 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.13 LAYER li1 ;
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.145 0.455 1.815 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER li1 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.3 5.205 6.61 5.875 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.06 LAYER li1 ;
  END CLK

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.64 5.6 7.81 6.235 ;
        RECT 5.305 6.235 7.81 6.405 ;
        RECT 5.305 5.525 5.475 6.235 ;
        RECT 5.145 4.885 5.475 5.525 ;
        RECT 7.64 5.535 8.485 5.6 ;
        RECT 8.3 5.205 8.89 5.43 ;
        RECT 7.64 5.43 8.89 5.535 ;
    END
    ANTENNAGATEAREA 0.598 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.191 LAYER li1 ;
  END SLEEPB

  PIN SETB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met1 ;
        RECT 2.14 2.705 15.365 2.845 ;
        RECT 14.715 2.845 15.365 2.92 ;
        RECT 14.715 2.69 15.365 2.705 ;
        RECT 2.14 2.845 2.795 2.92 ;
        RECT 8.235 2.845 8.885 2.92 ;
        RECT 2.14 2.69 2.795 2.705 ;
        RECT 8.235 2.69 8.885 2.705 ;
    END
    ANTENNAGATEAREA 0.378 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 9.3065 LAYER met1 ;
  END SETB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 16.8 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 16.8 6.905 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 16.8 3.575 ;
        RECT 2.975 3.075 6.145 3.085 ;
        RECT 11.85 2.985 13.33 3.085 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 3.715 16.73 3.985 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 13.04 3.285 13.21 3.455 ;
      RECT 12.645 3.075 12.815 3.245 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 6.575 12.805 6.745 ;
      RECT 12.285 3.075 12.455 3.245 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 6.575 12.325 6.745 ;
      RECT 11.915 3.03 12.085 3.2 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 6.575 11.845 6.745 ;
      RECT 11.54 3.785 11.71 3.955 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 6.575 11.365 6.745 ;
      RECT 11.18 3.785 11.35 3.955 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 6.575 10.885 6.745 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 6.155 3.785 6.325 3.955 ;
      RECT 5.265 3.785 5.435 3.955 ;
      RECT 10.235 6.575 10.405 6.745 ;
      RECT 5.915 3.105 6.085 3.275 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 6.575 9.925 6.745 ;
      RECT 9.615 3.245 9.785 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 6.575 9.445 6.745 ;
      RECT 9.255 3.18 9.425 3.35 ;
      RECT 8.895 3.18 9.065 3.35 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 6.575 8.965 6.745 ;
      RECT 8.655 2.72 8.825 2.89 ;
      RECT 8.535 3.18 8.705 3.35 ;
      RECT 8.295 2.72 8.465 2.89 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 6.575 8.485 6.745 ;
      RECT 8.255 3.765 8.425 3.935 ;
      RECT 8.175 3.18 8.345 3.35 ;
      RECT 7.895 3.765 8.065 3.935 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 6.575 8.005 6.745 ;
      RECT 7.815 3.18 7.985 3.35 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 7.455 3.18 7.625 3.35 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 6.575 7.525 6.745 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 6.575 7.045 6.745 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.555 3.105 5.725 3.275 ;
      RECT 6.395 6.575 6.565 6.745 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.195 3.105 5.365 3.275 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 4.835 3.105 5.005 3.275 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 4.475 3.105 4.645 3.275 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 4.115 3.105 4.285 3.275 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.755 3.105 3.925 3.275 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.395 3.105 3.565 3.275 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.105 3.205 3.275 ;
      RECT 3.035 6.575 3.205 6.745 ;
      RECT 2.56 2.72 2.73 2.89 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 2.2 2.72 2.37 2.89 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 16.475 6.575 16.645 6.745 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.995 6.575 16.165 6.745 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.515 6.575 15.685 6.745 ;
      RECT 15.155 3.295 15.325 3.465 ;
      RECT 15.135 2.72 15.305 2.89 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 6.575 15.205 6.745 ;
      RECT 14.795 3.295 14.965 3.465 ;
      RECT 14.775 2.72 14.945 2.89 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 6.575 14.725 6.745 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 6.575 14.245 6.745 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 6.575 13.765 6.745 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 6.575 13.285 6.745 ;
    LAYER li1 ;
      RECT 6.82 5.475 7.18 5.69 ;
      RECT 6.82 5.69 7.47 6.065 ;
      RECT 4.215 3.925 4.995 4.595 ;
      RECT 4.215 4.595 4.54 5.285 ;
      RECT 3.505 5.285 4.54 5.455 ;
      RECT 3.505 5.455 3.675 5.535 ;
      RECT 4.28 5.455 4.54 5.955 ;
      RECT 3.415 5.535 3.675 5.955 ;
      RECT 10.46 3.605 10.96 4.685 ;
      RECT 10.745 3.585 10.96 3.605 ;
      RECT 10.46 4.685 10.63 5.69 ;
      RECT 10.745 3.415 12.77 3.585 ;
      RECT 10.46 5.69 10.8 6.02 ;
      RECT 12.49 3.585 12.77 4.305 ;
      RECT 11.13 3.755 11.79 4.685 ;
      RECT 11.99 3.755 12.32 4.875 ;
      RECT 11.99 4.875 13.465 4.91 ;
      RECT 10.8 4.91 13.465 5.11 ;
      RECT 10.8 5.11 11.05 5.24 ;
      RECT 12.47 5.11 13.465 5.19 ;
      RECT 12.47 5.19 12.705 6.02 ;
      RECT 8.525 4.155 9.36 4.865 ;
      RECT 8.6 3.795 9.36 4.155 ;
      RECT 7.365 4.865 9.36 5.035 ;
      RECT 9.03 3.73 9.36 3.795 ;
      RECT 9.06 5.035 9.36 5.38 ;
      RECT 9.06 5.38 9.91 5.55 ;
      RECT 9.06 5.55 9.23 5.705 ;
      RECT 9.74 5.55 9.91 6.19 ;
      RECT 8.77 5.705 9.23 6.065 ;
      RECT 9.74 6.19 11.34 6.39 ;
      RECT 11.17 5.55 11.34 6.19 ;
      RECT 11.17 5.38 12.3 5.55 ;
      RECT 12.13 5.55 12.3 6.19 ;
      RECT 11.225 5.285 12.3 5.38 ;
      RECT 12.13 6.19 13.445 6.39 ;
      RECT 13.135 5.525 13.445 6.19 ;
      RECT 7.365 5.035 8.035 5.26 ;
      RECT 11.915 2.87 13.305 3.245 ;
      RECT 11.915 1.895 12.295 2.87 ;
      RECT 12.94 3.245 13.305 4.065 ;
      RECT 12.94 4.065 13.415 4.395 ;
      RECT 15.15 4.23 15.4 4.775 ;
      RECT 15.15 4.775 16.3 4.945 ;
      RECT 16.07 4.23 16.3 4.775 ;
      RECT 14.775 2.455 15.305 3.125 ;
      RECT 14.435 3.295 16.8 3.415 ;
      RECT 15.475 3.245 16.8 3.295 ;
      RECT 15.57 3.575 15.9 4.605 ;
      RECT 14.435 3.415 15.9 3.575 ;
      RECT 14.435 2.19 14.605 3.295 ;
      RECT 15.475 2.19 15.825 3.245 ;
      RECT 14.435 1.84 15.825 2.19 ;
      RECT 13.975 3.745 14.345 4.275 ;
      RECT 13.975 2.65 14.265 3.745 ;
      RECT 13.975 4.275 14.915 5.16 ;
      RECT 13.975 5.16 14.235 5.33 ;
      RECT 14.745 5.16 14.915 5.72 ;
      RECT 13.615 5.33 14.235 5.66 ;
      RECT 14.745 5.72 15.095 6.05 ;
      RECT 6.38 0.255 8.73 0.425 ;
      RECT 8.56 0.425 8.73 1.03 ;
      RECT 8.56 1.03 10.455 1.125 ;
      RECT 7.925 1.125 10.455 1.2 ;
      RECT 10.285 0.425 10.455 1.03 ;
      RECT 7.925 1.2 8.73 1.295 ;
      RECT 10.285 0.255 11.82 0.425 ;
      RECT 7.925 1.295 8.515 1.455 ;
      RECT 11.65 0.425 11.82 1.11 ;
      RECT 11.65 1.11 13.09 1.345 ;
      RECT 12.835 1.345 13.09 2.31 ;
      RECT 3.85 3.615 4.02 4.945 ;
      RECT 2.825 4.945 4.02 5.115 ;
      RECT 2.825 5.115 3.335 5.365 ;
      RECT 6.38 0.425 6.63 3.445 ;
      RECT 3.85 3.445 6.63 3.615 ;
      RECT 0 -0.085 16.8 0.085 ;
      RECT 0.965 0.085 1.3 1.06 ;
      RECT 2.93 0.085 3.25 1.015 ;
      RECT 4.56 0.085 4.81 0.975 ;
      RECT 5.88 0.085 6.21 0.955 ;
      RECT 9.21 0.085 10.115 0.86 ;
      RECT 11.99 0.085 15.825 0.285 ;
      RECT 11.99 0.285 12.645 0.94 ;
      RECT 14.405 0.285 15.825 1.07 ;
      RECT 0 6.575 16.8 6.745 ;
      RECT 8.01 6.265 9.57 6.575 ;
      RECT 11.51 5.72 11.96 6.575 ;
      RECT 14.28 6.22 16.285 6.575 ;
      RECT 8.01 5.77 8.6 6.265 ;
      RECT 9.4 5.72 9.57 6.265 ;
      RECT 14.28 5.83 14.575 6.22 ;
      RECT 15.955 5.72 16.285 6.22 ;
      RECT 14.405 5.33 14.575 5.83 ;
      RECT 1.1 6.28 4.11 6.575 ;
      RECT 4.73 5.68 5.06 6.575 ;
      RECT 2.05 5.625 2.315 6.28 ;
      RECT 2.915 5.625 3.245 6.28 ;
      RECT 3.845 5.625 4.11 6.28 ;
      RECT 1.1 5.605 1.395 6.28 ;
      RECT 4.98 0.645 5.6 0.975 ;
      RECT 3.975 1.32 4.225 1.815 ;
      RECT 3.975 1.145 5.15 1.32 ;
      RECT 4.85 1.32 5.1 2.655 ;
      RECT 4.98 0.975 5.15 1.145 ;
      RECT 3.585 0.975 3.805 1.985 ;
      RECT 3.45 0.255 4.1 0.975 ;
      RECT 3.585 1.985 4.14 2.205 ;
      RECT 3.91 2.205 4.14 2.655 ;
      RECT 2.495 1.185 3.415 1.855 ;
      RECT 2.495 0.65 2.76 1.185 ;
      RECT 2.495 1.855 2.76 2.34 ;
      RECT 1.97 0.975 2.19 1.99 ;
      RECT 1.675 0.255 2.325 0.975 ;
      RECT 1.515 1.99 2.19 2.175 ;
      RECT 1.515 2.175 1.785 2.66 ;
      RECT 0.625 1.615 1.8 1.82 ;
      RECT 1.55 1.145 1.8 1.615 ;
      RECT 0.625 0.975 0.795 1.615 ;
      RECT 0.625 1.82 0.845 2.66 ;
      RECT 0.095 0.645 0.795 0.975 ;
      RECT 7.575 1.71 9.615 1.88 ;
      RECT 7.575 1.185 7.755 1.71 ;
      RECT 8.28 1.88 8.49 2.345 ;
      RECT 9.345 1.88 9.615 2.335 ;
      RECT 7.305 0.955 7.755 1.185 ;
      RECT 7.305 0.595 8.39 0.955 ;
      RECT 10.585 1.59 10.895 2.38 ;
      RECT 10.045 1.54 10.895 1.59 ;
      RECT 9.065 1.37 10.895 1.54 ;
      RECT 10.625 0.625 10.895 1.37 ;
      RECT 11.145 1.725 11.46 3.025 ;
      RECT 11.145 1.515 12.665 1.725 ;
      RECT 10.225 3.025 11.46 3.245 ;
      RECT 12.465 1.725 12.665 2.48 ;
      RECT 11.145 0.595 11.48 1.515 ;
      RECT 10.225 3.245 10.575 3.435 ;
      RECT 12.465 2.48 13.805 2.7 ;
      RECT 13.26 1.67 13.805 2.48 ;
      RECT 13.475 2.7 13.805 3.68 ;
      RECT 13.26 1.24 15.825 1.67 ;
      RECT 13.26 0.755 13.97 1.24 ;
      RECT 2.895 3.275 3.265 4.775 ;
      RECT 2.895 3.24 6.21 3.275 ;
      RECT 2.93 2.855 6.21 3.24 ;
      RECT 2.93 2.025 3.28 2.855 ;
      RECT 4.315 2.835 6.21 2.855 ;
      RECT 5.27 2.015 6.21 2.835 ;
      RECT 4.315 1.985 4.68 2.835 ;
      RECT 2.14 2.61 2.76 2.94 ;
      RECT 1.59 3.84 1.99 4.64 ;
      RECT 0.895 3.585 1.99 3.84 ;
      RECT 1.59 4.64 2.655 4.84 ;
      RECT 1.59 4.84 1.88 5.955 ;
      RECT 2.485 4.84 2.655 5.535 ;
      RECT 2.485 5.535 2.745 5.955 ;
      RECT 0 3.245 1.345 3.415 ;
      RECT 0.095 2.84 1.345 3.245 ;
      RECT 1.015 1.99 1.345 2.84 ;
      RECT 0.16 3.415 0.52 4.84 ;
      RECT 0.095 2.02 0.455 2.84 ;
      RECT 0.69 4.17 0.93 5.255 ;
      RECT 0.235 5.255 0.93 5.955 ;
      RECT 7.365 3.09 9.81 3.535 ;
      RECT 9.53 3.535 9.81 4.685 ;
      RECT 9.005 2.855 9.81 3.09 ;
      RECT 9.005 2.505 10.385 2.855 ;
      RECT 9.005 2.345 9.175 2.505 ;
      RECT 10.045 1.99 10.385 2.505 ;
      RECT 8.66 2.05 9.175 2.345 ;
      RECT 8.245 2.54 8.835 2.92 ;
      RECT 7.965 3.985 8.355 4.695 ;
      RECT 7.89 3.705 8.43 3.985 ;
      RECT 5.235 3.955 5.475 4.715 ;
      RECT 5.235 3.785 6.355 3.955 ;
      RECT 6.145 3.955 6.355 4.695 ;
      RECT 6.525 4.23 6.695 4.865 ;
      RECT 6.525 4.06 6.97 4.23 ;
      RECT 6.8 2.895 6.97 4.06 ;
      RECT 6.8 2.225 7.13 2.895 ;
      RECT 5.645 4.865 6.695 5.035 ;
      RECT 5.645 4.125 5.975 4.865 ;
      RECT 5.92 5.035 6.13 6.01 ;
      RECT 7.465 4.155 7.795 4.525 ;
      RECT 7.465 3.795 7.72 4.155 ;
      RECT 7.01 4.525 7.795 4.695 ;
      RECT 7.01 4.695 7.18 5.475 ;
  END
END scs8ls_lpflow_srsdfstp2_1

MACRO scs8ls_lpflow_srsdfrtp2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 17.28 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.5 1.125 6.085 1.44 ;
        RECT 5.5 1.44 5.725 1.795 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.183 LAYER li1 ;
  END SCD

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.725 0.37 17.155 3.015 ;
    END
    ANTENNADIFFAREA 0.5097 ;
    ANTENNAPARTIALMETALSIDEAREA 0.547 LAYER li1 ;
  END Q

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.49 5.035 2.08 5.455 ;
    END
    ANTENNAGATEAREA 0.318 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.134 LAYER li1 ;
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.095 0.425 1.765 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.058 LAYER li1 ;
  END D

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.68 4.895 7.195 5.515 ;
    END
    ANTENNAGATEAREA 0.159 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.091 LAYER li1 ;
  END CLK

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.15 5.205 9.85 5.38 ;
        RECT 8.615 5.38 9.85 5.535 ;
        RECT 8.615 5.535 9.32 5.55 ;
        RECT 8.615 5.55 8.785 6.235 ;
        RECT 7.225 6.235 8.785 6.405 ;
        RECT 7.225 6.205 7.595 6.235 ;
        RECT 7.425 5.265 7.595 6.205 ;
        RECT 7.425 4.935 7.74 5.265 ;
    END
    ANTENNAGATEAREA 0.598 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.986 LAYER li1 ;
  END SLEEPB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 17.28 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 17.28 6.905 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 17.28 3.575 ;
        RECT 6.38 2.985 8.11 3.085 ;
        RECT 10.405 2.985 15.03 3.085 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 3.715 17.21 3.985 ;
    END
  END kapwr

  PIN RESETB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met1 ;
        RECT 2.535 2.705 15.83 2.845 ;
        RECT 15.17 2.845 15.83 2.935 ;
        RECT 15.515 2.69 15.83 2.705 ;
        RECT 2.535 2.845 3.215 2.935 ;
        RECT 8.45 2.845 9.1 2.92 ;
        RECT 2.535 2.69 3.215 2.705 ;
        RECT 8.45 2.69 9.1 2.705 ;
    END
    ANTENNAGATEAREA 0.378 LAYER met1 ;
    ANTENNAPARTIALMETALSIDEAREA 9.3765 LAYER met1 ;
  END RESETB

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 6.575 15.205 6.745 ;
      RECT 14.8 3.015 14.97 3.185 ;
      RECT 14.8 3.375 14.97 3.545 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 6.575 14.725 6.745 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 6.575 14.245 6.745 ;
      RECT 13.95 3.015 14.12 3.185 ;
      RECT 13.95 3.375 14.12 3.545 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 6.575 13.765 6.745 ;
      RECT 13.59 3.015 13.76 3.185 ;
      RECT 13.23 3.015 13.4 3.185 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 6.575 13.285 6.745 ;
      RECT 12.87 3.015 13.04 3.185 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 6.575 12.805 6.745 ;
      RECT 12.51 3.015 12.68 3.185 ;
      RECT 12.5 3.785 12.67 3.955 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 6.575 12.325 6.745 ;
      RECT 12.14 3.785 12.31 3.955 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 6.575 11.845 6.745 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 6.575 11.365 6.745 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 6.575 10.885 6.745 ;
      RECT 10.51 3.375 10.68 3.545 ;
      RECT 10.465 3.015 10.635 3.185 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 6.575 10.405 6.745 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 6.575 9.925 6.745 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 6.575 9.445 6.745 ;
      RECT 9.215 3.765 9.385 3.935 ;
      RECT 8.87 2.72 9.04 2.89 ;
      RECT 8.855 3.765 9.025 3.935 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 6.575 8.965 6.745 ;
      RECT 8.51 2.72 8.68 2.89 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 6.575 8.485 6.745 ;
      RECT 8.04 3.785 8.21 3.955 ;
      RECT 7.88 3.105 8.05 3.275 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 6.575 8.005 6.745 ;
      RECT 7.68 3.785 7.85 3.955 ;
      RECT 7.52 3.105 7.69 3.275 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 6.575 7.525 6.745 ;
      RECT 7.16 3.105 7.33 3.275 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 6.575 7.045 6.745 ;
      RECT 6.8 3.105 6.97 3.275 ;
      RECT 6.795 3.785 6.965 3.955 ;
      RECT 6.44 3.015 6.61 3.185 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 6.575 6.565 6.745 ;
      RECT 6.315 3.375 6.485 3.545 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 5.475 3.245 5.645 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 5.105 3.245 5.275 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 16.995 3.245 17.165 3.415 ;
      RECT 16.955 -0.085 17.125 0.085 ;
      RECT 16.955 6.575 17.125 6.745 ;
      RECT 16.635 3.245 16.805 3.415 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 16.475 6.575 16.645 6.745 ;
      RECT 16.275 3.295 16.445 3.465 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 6.575 16.165 6.745 ;
      RECT 15.915 3.295 16.085 3.465 ;
      RECT 15.6 2.735 15.77 2.905 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 4.525 3.245 4.695 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 4.155 3.245 4.325 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 3.785 3.245 3.955 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 3.415 3.245 3.585 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 6.575 3.205 6.745 ;
      RECT 2.985 2.735 3.155 2.905 ;
      RECT 2.595 2.735 2.765 2.905 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 1.26 3.245 1.43 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 0.89 3.245 1.06 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 0.525 3.245 0.695 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 6.575 15.685 6.745 ;
      RECT 15.24 2.735 15.41 2.905 ;
    LAYER li1 ;
      RECT 3.355 2.79 5.725 3.415 ;
      RECT 3.355 2.525 3.825 2.79 ;
      RECT 5.385 1.97 5.725 2.79 ;
      RECT 4.475 1.935 4.805 2.79 ;
      RECT 3.115 2.315 3.825 2.525 ;
      RECT 3.115 1.925 3.445 2.315 ;
      RECT 4.77 4.17 5.54 4.595 ;
      RECT 5.21 3.925 5.54 4.17 ;
      RECT 4.77 4.595 5.09 5.43 ;
      RECT 4.005 5.43 5.13 5.6 ;
      RECT 4.005 5.6 4.195 5.995 ;
      RECT 4.88 5.6 5.13 5.955 ;
      RECT 2.565 2.695 3.185 3.025 ;
      RECT 9.485 4.155 9.815 4.865 ;
      RECT 9.56 4.11 9.815 4.155 ;
      RECT 8.81 4.865 10.19 4.955 ;
      RECT 9.56 3.795 10.32 4.11 ;
      RECT 8.31 4.955 10.19 5.035 ;
      RECT 9.99 3.52 10.32 3.795 ;
      RECT 10.02 5.035 10.19 5.38 ;
      RECT 10.02 5.38 11.22 5.55 ;
      RECT 10.02 5.55 10.19 5.735 ;
      RECT 11.05 5.55 11.22 6.22 ;
      RECT 9.825 5.735 10.19 6.065 ;
      RECT 11.05 6.22 12.3 6.39 ;
      RECT 12.13 5.55 12.3 6.22 ;
      RECT 12.13 5.38 13.26 5.55 ;
      RECT 13.09 5.55 13.26 6.22 ;
      RECT 12.345 5.285 12.675 5.38 ;
      RECT 13.09 6.22 14.425 6.39 ;
      RECT 14.095 5.865 14.425 6.22 ;
      RECT 14.095 5.525 14.405 5.865 ;
      RECT 8.31 5.035 8.98 5.21 ;
      RECT 8.955 3.985 9.285 4.695 ;
      RECT 8.85 3.705 9.39 3.985 ;
      RECT 8.41 2.655 9.14 2.93 ;
      RECT 8.41 1.935 9.08 2.655 ;
      RECT 8.425 4.155 8.755 4.615 ;
      RECT 8.425 3.795 8.68 4.155 ;
      RECT 7.97 4.615 8.755 4.695 ;
      RECT 7.97 4.695 8.595 4.785 ;
      RECT 7.97 4.785 8.14 5.475 ;
      RECT 7.765 5.475 8.14 5.735 ;
      RECT 7.765 5.735 8.445 6.065 ;
      RECT 7.635 3.785 8.255 4.445 ;
      RECT 6.275 3.275 6.525 4.385 ;
      RECT 6.275 3.085 8.15 3.275 ;
      RECT 6.275 1.95 6.69 3.085 ;
      RECT 7.855 1.93 8.15 3.085 ;
      RECT 6.715 3.705 7.045 4.385 ;
      RECT 12.45 2.955 14.17 3.245 ;
      RECT 12.45 1.945 13.03 2.955 ;
      RECT 13.9 3.245 14.17 4.165 ;
      RECT 12.745 1.825 13.03 1.945 ;
      RECT 13.9 4.165 14.455 4.445 ;
      RECT 11.42 3.585 11.795 4.685 ;
      RECT 11.42 3.415 13.73 3.585 ;
      RECT 11.42 4.685 11.59 5.72 ;
      RECT 13.45 3.585 13.73 4.305 ;
      RECT 11.42 5.72 11.76 6.05 ;
      RECT 12.42 3.985 12.75 4.685 ;
      RECT 12.09 3.755 12.75 3.985 ;
      RECT 10.49 3.4 10.78 4.685 ;
      RECT 10.49 3.35 10.695 3.4 ;
      RECT 10.405 2.73 10.695 3.35 ;
      RECT 10.405 1.97 10.77 2.73 ;
      RECT 12.95 3.755 13.28 4.94 ;
      RECT 11.76 4.94 14.855 5.11 ;
      RECT 11.76 5.11 12.01 5.24 ;
      RECT 13.45 5.11 13.7 6.05 ;
      RECT 11.76 4.91 12.01 4.94 ;
      RECT 14.265 5.11 14.855 5.16 ;
      RECT 14.265 4.83 14.855 4.94 ;
      RECT 15.18 2.935 15.43 3.4 ;
      RECT 15.18 2.705 15.83 2.935 ;
      RECT 14.76 2.25 15.01 3.575 ;
      RECT 14.505 1.92 15.01 2.25 ;
      RECT 15.025 4.995 16.955 5.165 ;
      RECT 16.625 5.165 16.955 6.05 ;
      RECT 16.45 4.275 16.78 4.995 ;
      RECT 14.66 4.045 15.265 4.215 ;
      RECT 14.66 3.995 14.91 4.045 ;
      RECT 15.025 4.215 15.265 4.995 ;
      RECT 14.34 3.745 14.91 3.995 ;
      RECT 14.34 2.88 14.59 3.745 ;
      RECT 15.025 5.165 15.195 5.33 ;
      RECT 14.575 5.33 15.195 5.5 ;
      RECT 14.575 5.5 14.825 5.685 ;
      RECT 15.6 3.415 16.75 4.075 ;
      RECT 15.6 3.295 17.28 3.415 ;
      RECT 16.265 3.245 17.28 3.295 ;
      RECT 15.6 4.075 15.93 4.605 ;
      RECT 16.265 1.855 16.515 3.245 ;
      RECT 0 6.575 17.28 6.745 ;
      RECT 8.955 5.72 9.285 6.575 ;
      RECT 10.36 5.72 10.75 6.575 ;
      RECT 12.5 5.72 12.89 6.575 ;
      RECT 15.365 5.72 16.085 6.575 ;
      RECT 15.365 5.355 15.615 5.72 ;
      RECT 1.51 5.625 1.775 6.575 ;
      RECT 2.64 5.77 2.97 6.575 ;
      RECT 4.37 5.77 4.7 6.575 ;
      RECT 5.84 5.67 6.17 6.575 ;
      RECT 3.505 5.625 3.835 6.575 ;
      RECT 0 -0.085 17.28 0.085 ;
      RECT 1.03 0.085 1.36 0.97 ;
      RECT 3.085 0.085 3.405 0.99 ;
      RECT 4.615 0.085 4.935 1 ;
      RECT 6.02 0.085 6.35 0.86 ;
      RECT 8.115 0.085 8.325 0.94 ;
      RECT 10.415 0.085 11.825 0.97 ;
      RECT 14.945 0.085 15.195 1.05 ;
      RECT 16.255 0.085 16.555 1.07 ;
      RECT 1.74 0.57 2.39 0.895 ;
      RECT 2.115 0.895 2.39 0.925 ;
      RECT 2.14 0.255 2.39 0.57 ;
      RECT 2.115 0.925 2.325 1.935 ;
      RECT 1.62 1.935 2.325 2.145 ;
      RECT 1.62 2.145 1.91 2.605 ;
      RECT 0.69 1.35 0.91 2.605 ;
      RECT 0.69 1.18 1.945 1.35 ;
      RECT 1.615 1.35 1.945 1.735 ;
      RECT 1.615 1.125 1.945 1.18 ;
      RECT 0.69 0.925 0.86 1.18 ;
      RECT 0.16 0.595 0.86 0.925 ;
      RECT 5.105 0.625 5.805 0.955 ;
      RECT 4.02 1.63 4.35 1.735 ;
      RECT 4.02 1.415 5.33 1.63 ;
      RECT 4.975 1.63 5.215 2.605 ;
      RECT 4.02 1.125 4.35 1.415 ;
      RECT 5.105 0.955 5.33 1.415 ;
      RECT 3.64 0.925 3.85 1.935 ;
      RECT 3.575 0.6 4.225 0.925 ;
      RECT 3.64 1.935 4.265 2.145 ;
      RECT 3.575 0.255 3.825 0.6 ;
      RECT 4.055 2.145 4.265 2.605 ;
      RECT 2.495 1.095 2.915 1.825 ;
      RECT 2.645 0.64 2.915 1.095 ;
      RECT 2.66 1.825 2.915 2.34 ;
      RECT 8.495 0.255 10.245 0.425 ;
      RECT 10.075 0.425 10.245 1.15 ;
      RECT 10.075 1.15 12.165 1.32 ;
      RECT 10.075 1.32 10.925 1.46 ;
      RECT 11.995 0.425 12.165 1.15 ;
      RECT 11.995 0.255 13.445 0.425 ;
      RECT 13.275 0.425 13.445 0.465 ;
      RECT 13.275 0.465 13.555 1.135 ;
      RECT 5.895 1.61 6.69 1.78 ;
      RECT 6.52 0.425 6.69 1.61 ;
      RECT 5.895 1.78 6.105 3.585 ;
      RECT 4.035 3.585 6.105 3.755 ;
      RECT 5.775 3.755 6.105 4.155 ;
      RECT 5.71 4.155 6.105 4.365 ;
      RECT 5.71 4.365 5.92 5.29 ;
      RECT 5.46 5.29 5.92 5.5 ;
      RECT 5.46 5.5 5.67 6.02 ;
      RECT 4.035 3.755 4.205 4.945 ;
      RECT 3.335 4.945 4.205 5.115 ;
      RECT 3.335 5.115 4.005 5.26 ;
      RECT 6.52 0.255 7.945 0.425 ;
      RECT 7.775 0.425 7.945 1.12 ;
      RECT 7.775 1.12 8.665 1.29 ;
      RECT 8.495 0.425 8.665 1.12 ;
      RECT 9.38 1.305 9.55 1.93 ;
      RECT 9.19 0.94 9.55 1.305 ;
      RECT 9.25 1.93 9.55 2.26 ;
      RECT 8.835 0.595 9.905 0.94 ;
      RECT 7.395 1.475 9.21 1.665 ;
      RECT 7.395 0.61 7.605 1.475 ;
      RECT 7.395 1.665 7.655 2.26 ;
      RECT 8.54 1.665 9.21 1.725 ;
      RECT 6.86 0.61 7.1 2.645 ;
      RECT 6.86 2.645 7.685 2.895 ;
      RECT 9.98 1.63 11.22 1.8 ;
      RECT 9.98 1.8 10.15 3.135 ;
      RECT 10.94 1.8 11.22 2.69 ;
      RECT 8.51 3.135 10.15 3.305 ;
      RECT 6.34 5.685 7.255 6.015 ;
      RECT 6.18 4.725 6.51 5.21 ;
      RECT 6.34 5.21 6.51 5.685 ;
      RECT 7.295 3.615 7.465 3.705 ;
      RECT 7.215 3.705 7.465 4.555 ;
      RECT 6.18 4.555 7.465 4.725 ;
      RECT 8.51 3.305 8.68 3.445 ;
      RECT 7.295 3.445 8.68 3.615 ;
      RECT 11.85 1.49 12.575 1.775 ;
      RECT 12.335 1.475 12.575 1.49 ;
      RECT 11.85 1.775 12.18 2.9 ;
      RECT 12.335 1.305 13.975 1.475 ;
      RECT 10.865 2.9 12.18 3.07 ;
      RECT 12.335 0.625 12.575 1.305 ;
      RECT 13.675 1.475 13.975 1.56 ;
      RECT 13.725 0.72 13.975 1.305 ;
      RECT 10.865 3.07 11.455 3.23 ;
      RECT 13.675 1.56 16.555 1.625 ;
      RECT 13.675 1.625 16.095 1.73 ;
      RECT 15.925 1.455 16.555 1.56 ;
      RECT 13.675 1.73 13.965 2.295 ;
      RECT 15.375 1.73 15.665 2.295 ;
      RECT 15.965 1.295 16.555 1.455 ;
      RECT 14.475 1.22 15.625 1.39 ;
      RECT 14.475 0.72 14.775 1.22 ;
      RECT 15.365 0.72 15.625 1.22 ;
      RECT 0.505 4.11 0.87 4.84 ;
      RECT 0.505 3.415 0.725 4.11 ;
      RECT 0 3.245 1.46 3.415 ;
      RECT 0.22 2.79 1.46 3.245 ;
      RECT 0.22 2.785 1.41 2.79 ;
      RECT 0.22 1.935 0.5 2.785 ;
      RECT 1.08 1.935 1.41 2.785 ;
      RECT 1.08 4.17 1.32 5.255 ;
      RECT 0.6 5.255 1.32 5.925 ;
      RECT 1.08 5.925 1.32 5.955 ;
      RECT 0.925 3.585 2.61 3.84 ;
      RECT 2.25 3.84 2.61 4.845 ;
      RECT 2.25 4.845 2.46 5.43 ;
      RECT 2.25 5.43 3.335 5.6 ;
      RECT 2.25 5.6 2.46 5.955 ;
      RECT 3.145 5.6 3.335 5.995 ;
      RECT 3.505 3.415 3.835 4.775 ;
  END
END scs8ls_lpflow_srsdfrtp2_1

MACRO scs8ls_lpflow_lsbuf_lh_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.6 0.8 7.085 1.82 ;
        RECT 6.565 1.82 7.085 2.16 ;
        RECT 6.6 0.35 6.82 0.8 ;
        RECT 6.565 2.16 6.76 2.98 ;
    END
    ANTENNADIFFAREA 0.5041 ;
    ANTENNAPARTIALMETALSIDEAREA 0.358 LAYER li1 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045 2.23 1.325 2.53 ;
        RECT 1.045 1.9 1.665 2.23 ;
    END
    ANTENNAGATEAREA 0.675 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.114 LAYER li1 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
    END
  END vpwr

  PIN lowlvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 7.13 2.945 ;
    END
  END lowlvpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 5.585 1.63 5.795 2.98 ;
      RECT 5.585 1.3 6.43 1.63 ;
      RECT 5.64 0.35 5.855 1.3 ;
      RECT 0 -0.085 7.2 0.085 ;
      RECT 6.1 0.085 6.43 1.13 ;
      RECT 3.485 0.085 3.76 1.05 ;
      RECT 4.29 0.085 4.62 1.05 ;
      RECT 5.15 0.085 5.47 1.13 ;
      RECT 2.305 0.085 2.635 1.05 ;
      RECT 0.585 0.085 0.915 1.13 ;
      RECT 1.445 0.085 1.775 1.05 ;
      RECT 0 3.245 7.2 3.415 ;
      RECT 5.075 1.82 5.405 3.245 ;
      RECT 6.045 1.82 6.375 3.245 ;
      RECT 3.11 1.9 3.35 3.245 ;
      RECT 0.545 2.7 1.555 2.97 ;
      RECT 0.545 1.9 0.875 2.7 ;
      RECT 3.86 1.39 4.03 2.735 ;
      RECT 3.11 1.22 4.98 1.39 ;
      RECT 3.11 0.72 3.28 1.22 ;
      RECT 3.93 0.35 4.12 1.22 ;
      RECT 4.285 1.39 4.905 1.78 ;
      RECT 4.79 0.35 4.98 1.22 ;
      RECT 3.52 2.905 4.56 3.075 ;
      RECT 4.23 2.29 4.56 2.905 ;
      RECT 3.52 1.73 3.69 2.905 ;
      RECT 2.7 1.56 3.69 1.73 ;
      RECT 2.7 1.73 2.94 3.005 ;
      RECT 2.7 1.39 2.94 1.56 ;
      RECT 1.085 1.22 2.94 1.39 ;
      RECT 1.085 0.35 1.275 1.22 ;
      RECT 1.945 0.35 2.135 1.22 ;
      RECT 0.135 1.56 2.53 1.73 ;
      RECT 2.2 1.73 2.53 2.215 ;
      RECT 0.135 1.73 0.375 2.98 ;
      RECT 0.135 0.735 0.375 1.56 ;
    LAYER mcon ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.625 2.715 0.795 2.885 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 1.345 2.725 1.515 2.895 ;
      RECT 0.985 2.725 1.155 2.895 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
  END
END scs8ls_lpflow_lsbuf_lh_1

MACRO scs8ls_lpflow_lsbuf_lh_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.68 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845 0.35 7.075 2.98 ;
    END
    ANTENNADIFFAREA 0.5432 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3 LAYER li1 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045 2.23 1.325 2.53 ;
        RECT 1.045 1.9 1.665 2.23 ;
    END
    ANTENNAGATEAREA 0.675 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.114 LAYER li1 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.68 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.68 3.575 ;
    END
  END vpwr

  PIN lowlvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 7.61 2.945 ;
    END
  END lowlvpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 5.585 1.63 5.795 2.98 ;
      RECT 5.585 1.3 6.675 1.63 ;
      RECT 5.64 0.35 5.855 1.3 ;
      RECT 0 -0.085 7.68 0.085 ;
      RECT 7.245 0.085 7.555 1.13 ;
      RECT 6.365 0.085 6.675 1.13 ;
      RECT 3.485 0.085 3.76 1.05 ;
      RECT 4.29 0.085 4.62 1.05 ;
      RECT 5.15 0.085 5.47 1.13 ;
      RECT 2.305 0.085 2.635 1.05 ;
      RECT 0.585 0.085 0.915 1.13 ;
      RECT 1.445 0.085 1.775 1.05 ;
      RECT 7.245 1.82 7.575 3.245 ;
      RECT 0 3.245 7.68 3.415 ;
      RECT 5.075 1.82 5.405 3.245 ;
      RECT 6.345 1.82 6.675 3.245 ;
      RECT 3.11 1.9 3.35 3.245 ;
      RECT 0.545 2.7 1.555 2.97 ;
      RECT 0.545 1.9 0.875 2.7 ;
      RECT 3.86 1.39 4.03 2.735 ;
      RECT 3.11 1.22 4.98 1.39 ;
      RECT 3.11 0.72 3.28 1.22 ;
      RECT 3.93 0.35 4.12 1.22 ;
      RECT 4.285 1.39 4.905 1.78 ;
      RECT 4.79 0.35 4.98 1.22 ;
      RECT 3.52 2.905 4.56 3.075 ;
      RECT 4.23 2.29 4.56 2.905 ;
      RECT 3.52 1.73 3.69 2.905 ;
      RECT 2.7 1.56 3.69 1.73 ;
      RECT 2.7 1.73 2.94 3.005 ;
      RECT 2.7 1.39 2.94 1.56 ;
      RECT 1.085 1.22 2.94 1.39 ;
      RECT 1.085 0.35 1.275 1.22 ;
      RECT 1.945 0.35 2.135 1.22 ;
      RECT 0.135 1.56 2.53 1.73 ;
      RECT 2.2 1.73 2.53 2.215 ;
      RECT 0.135 1.73 0.375 2.98 ;
      RECT 0.135 0.735 0.375 1.56 ;
    LAYER mcon ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.625 2.715 0.795 2.885 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 1.345 2.725 1.515 2.895 ;
      RECT 0.985 2.725 1.155 2.895 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
  END
END scs8ls_lpflow_lsbuf_lh_2

MACRO scs8ls_lpflow_lsbuf_lh_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805 0.35 8.035 1.365 ;
        RECT 6.905 1.365 8.035 1.595 ;
        RECT 6.905 1.595 7.135 2.98 ;
        RECT 7.805 1.595 8.035 2.98 ;
        RECT 6.945 0.35 7.175 1.365 ;
    END
    ANTENNADIFFAREA 1.0864 ;
    ANTENNAPARTIALMETALSIDEAREA 1.096 LAYER li1 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045 2.23 1.325 2.53 ;
        RECT 1.045 1.9 1.665 2.23 ;
    END
    ANTENNAGATEAREA 0.675 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.114 LAYER li1 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN lowlvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 8.57 2.945 ;
    END
  END lowlvpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 8.205 1.82 8.535 3.245 ;
      RECT 6.405 1.82 6.735 3.245 ;
      RECT 5.075 1.82 5.405 3.245 ;
      RECT 3.11 1.9 3.35 3.245 ;
      RECT 7.305 1.82 7.635 3.245 ;
      RECT 5.585 1.63 5.795 2.98 ;
      RECT 5.585 1.3 6.735 1.63 ;
      RECT 5.64 0.35 5.855 1.3 ;
      RECT 8.205 0.085 8.515 1.13 ;
      RECT 0 -0.085 8.64 0.085 ;
      RECT 6.485 0.085 6.775 1.13 ;
      RECT 3.485 0.085 3.76 1.05 ;
      RECT 4.29 0.085 4.62 1.05 ;
      RECT 5.15 0.085 5.47 1.13 ;
      RECT 2.305 0.085 2.635 1.05 ;
      RECT 0.585 0.085 0.915 1.13 ;
      RECT 1.445 0.085 1.775 1.05 ;
      RECT 7.345 0.085 7.635 1.13 ;
      RECT 0.545 2.7 1.555 2.97 ;
      RECT 0.545 1.9 0.875 2.7 ;
      RECT 3.86 1.39 4.03 2.735 ;
      RECT 3.11 1.22 4.98 1.39 ;
      RECT 3.11 0.72 3.28 1.22 ;
      RECT 3.93 0.35 4.12 1.22 ;
      RECT 4.285 1.39 4.905 1.78 ;
      RECT 4.79 0.35 4.98 1.22 ;
      RECT 3.52 2.905 4.56 3.075 ;
      RECT 4.23 2.29 4.56 2.905 ;
      RECT 3.52 1.73 3.69 2.905 ;
      RECT 2.7 1.56 3.69 1.73 ;
      RECT 2.7 1.73 2.94 3.005 ;
      RECT 2.7 1.39 2.94 1.56 ;
      RECT 1.085 1.22 2.94 1.39 ;
      RECT 1.085 0.35 1.275 1.22 ;
      RECT 1.945 0.35 2.135 1.22 ;
      RECT 0.135 1.56 2.53 1.73 ;
      RECT 2.2 1.73 2.53 2.215 ;
      RECT 0.135 1.73 0.375 2.98 ;
      RECT 0.135 0.735 0.375 1.56 ;
    LAYER mcon ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 1.345 2.725 1.515 2.895 ;
      RECT 0.985 2.725 1.155 2.895 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.625 2.715 0.795 2.885 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
  END
END scs8ls_lpflow_lsbuf_lh_4

MACRO scs8ls_lpflow_lsbuf_lh_isowell_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.24 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.36 1.55 5.635 2.98 ;
        RECT 5.335 0.35 5.635 1.55 ;
    END
    ANTENNADIFFAREA 0.5041 ;
    ANTENNAPARTIALMETALSIDEAREA 0.45 LAYER li1 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.83 3.29 2.15 ;
        RECT 2.97 1.56 3.63 1.83 ;
        RECT 2.97 1.5 3.445 1.56 ;
    END
    ANTENNAGATEAREA 0.675 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER li1 ;
  END A

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
    END
  END vpwr

  PIN lowlvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 6.17 2.945 ;
    END
  END lowlvpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 6.24 6.905 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.615 1.22 4.665 1.39 ;
      RECT 3.615 0.35 3.805 1.22 ;
      RECT 4.475 0.35 4.665 1.22 ;
      RECT 3.68 3.185 3.85 4.235 ;
      RECT 3.68 3.015 4.19 3.185 ;
      RECT 4.02 1.39 4.19 3.015 ;
      RECT 4.39 4.405 4.72 4.84 ;
      RECT 3.68 4.235 4.72 4.405 ;
      RECT 4.39 3.695 4.72 4.235 ;
      RECT 4.89 3.245 6.24 3.415 ;
      RECT 4.89 1.82 5.12 3.245 ;
      RECT 4.89 3.415 5.12 4.84 ;
      RECT 3.145 5.19 5.19 5.36 ;
      RECT 4.6 5.01 5.19 5.19 ;
      RECT 4.005 5.36 4.195 6.31 ;
      RECT 3.145 5.36 3.335 6.31 ;
      RECT 5.205 5.72 5.55 6.31 ;
      RECT 5.205 5.53 5.865 5.72 ;
      RECT 5.36 5.05 5.865 5.53 ;
      RECT 5.36 3.68 5.55 5.05 ;
      RECT 3.06 4.77 3.73 5.02 ;
      RECT 3.06 2.98 3.3 4.77 ;
      RECT 2.56 2.74 3.3 2.98 ;
      RECT 2.56 0.735 2.8 2.74 ;
      RECT 0 3.245 1.89 3.415 ;
      RECT 4.365 5.53 5.035 6.575 ;
      RECT 0 6.575 6.24 6.745 ;
      RECT 3.505 5.53 3.835 6.575 ;
      RECT 2.645 5.53 2.975 6.575 ;
      RECT 4.02 3.525 4.19 4.065 ;
      RECT 4.02 3.355 4.64 3.525 ;
      RECT 4.47 1.82 4.64 3.355 ;
      RECT 2.06 3.27 2.81 3.94 ;
      RECT 2.06 2.945 2.39 3.27 ;
      RECT 1.38 2.675 2.39 2.945 ;
      RECT 2.06 1.9 2.39 2.675 ;
      RECT 0 -0.085 6.24 0.085 ;
      RECT 3.115 0.085 3.445 1.13 ;
      RECT 3.975 0.085 4.305 1.05 ;
      RECT 4.835 0.085 5.165 1.13 ;
      RECT 2.02 0.085 2.35 1.13 ;
    LAYER mcon ;
      RECT 1.78 2.725 1.95 2.895 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 3.035 6.575 3.205 6.745 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.14 2.715 2.31 2.885 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 1.42 2.725 1.59 2.895 ;
  END
END scs8ls_lpflow_lsbuf_lh_isowell_1

MACRO scs8ls_lpflow_lsbuf_lh_isowell_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.24 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.355 1.3 5.685 2.98 ;
        RECT 5.355 0.35 5.59 1.3 ;
    END
    ANTENNADIFFAREA 0.5432 ;
    ANTENNAPARTIALMETALSIDEAREA 0.456 LAYER li1 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.83 3.29 2.15 ;
        RECT 2.97 1.56 3.63 1.83 ;
        RECT 2.97 1.5 3.445 1.56 ;
    END
    ANTENNAGATEAREA 0.675 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER li1 ;
  END A

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
    END
  END vpwr

  PIN lowlvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 6.17 2.945 ;
    END
  END lowlvpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 6.24 6.905 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 3.615 1.22 4.665 1.39 ;
      RECT 3.615 0.35 3.805 1.22 ;
      RECT 4.475 0.35 4.665 1.22 ;
      RECT 3.68 3.185 3.85 4.235 ;
      RECT 3.68 3.015 4.19 3.185 ;
      RECT 4.02 1.39 4.19 3.015 ;
      RECT 4.39 4.405 4.72 4.84 ;
      RECT 3.68 4.235 4.72 4.405 ;
      RECT 4.39 3.695 4.72 4.235 ;
      RECT 5.855 1.82 6.085 3.245 ;
      RECT 4.89 3.245 6.24 3.415 ;
      RECT 4.89 1.82 5.12 3.245 ;
      RECT 4.89 3.415 5.12 4.84 ;
      RECT 5.76 0.085 6.09 1.13 ;
      RECT 0 -0.085 6.24 0.085 ;
      RECT 3.115 0.085 3.445 1.13 ;
      RECT 3.975 0.085 4.305 1.05 ;
      RECT 4.835 0.085 5.165 1.13 ;
      RECT 2.02 0.085 2.35 1.13 ;
      RECT 3.145 5.19 5.19 5.36 ;
      RECT 4.6 5.01 5.19 5.19 ;
      RECT 4.005 5.36 4.195 6.31 ;
      RECT 3.145 5.36 3.335 6.31 ;
      RECT 5.205 5.72 5.55 6.31 ;
      RECT 5.205 5.53 5.865 5.72 ;
      RECT 5.36 5.05 5.865 5.53 ;
      RECT 5.36 3.68 5.55 5.05 ;
      RECT 3.06 4.77 3.73 5.02 ;
      RECT 3.06 2.98 3.3 4.77 ;
      RECT 2.56 2.74 3.3 2.98 ;
      RECT 2.56 0.735 2.8 2.74 ;
      RECT 0 3.245 1.89 3.415 ;
      RECT 4.365 5.53 5.035 6.575 ;
      RECT 0 6.575 6.24 6.745 ;
      RECT 3.505 5.53 3.835 6.575 ;
      RECT 2.645 5.53 2.975 6.575 ;
      RECT 4.02 3.525 4.19 4.065 ;
      RECT 4.02 3.355 4.64 3.525 ;
      RECT 4.47 1.82 4.64 3.355 ;
      RECT 2.06 3.27 2.81 3.94 ;
      RECT 2.06 2.945 2.39 3.27 ;
      RECT 1.38 2.675 2.39 2.945 ;
      RECT 2.06 1.9 2.39 2.675 ;
    LAYER mcon ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 1.42 2.725 1.59 2.895 ;
      RECT 1.78 2.725 1.95 2.895 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 3.035 6.575 3.205 6.745 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.14 2.715 2.31 2.885 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
  END
END scs8ls_lpflow_lsbuf_lh_isowell_2

MACRO scs8ls_lpflow_lsbuf_lh_isowell_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 6.66 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 1.59 6.595 2.98 ;
        RECT 5.465 1.36 6.595 1.59 ;
        RECT 5.465 1.59 5.695 2.98 ;
        RECT 5.465 0.35 5.695 1.36 ;
        RECT 6.365 0.35 6.595 1.36 ;
    END
    ANTENNADIFFAREA 1.0864 ;
    ANTENNAPARTIALMETALSIDEAREA 1.096 LAYER li1 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.83 3.29 2.15 ;
        RECT 2.97 1.56 3.63 1.83 ;
        RECT 2.97 1.5 3.445 1.56 ;
    END
    ANTENNAGATEAREA 0.675 LAYER li1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER li1 ;
  END A

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 7.2 3.575 ;
    END
  END vpwr

  PIN lowlvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 7.13 2.945 ;
    END
  END lowlvpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 7.2 0.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 6.415 7.2 6.905 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.645 5.53 2.975 6.575 ;
      RECT 0 6.575 7.2 6.745 ;
      RECT 4.365 5.53 5.035 6.575 ;
      RECT 3.505 5.53 3.835 6.575 ;
      RECT 4.02 3.525 4.19 4.065 ;
      RECT 4.02 3.355 4.64 3.525 ;
      RECT 4.47 1.82 4.64 3.355 ;
      RECT 2.06 3.27 2.81 3.94 ;
      RECT 2.06 2.945 2.39 3.27 ;
      RECT 1.38 2.675 2.39 2.945 ;
      RECT 2.06 1.9 2.39 2.675 ;
      RECT 4.89 3.245 7.2 3.415 ;
      RECT 6.765 1.82 7.095 3.245 ;
      RECT 4.89 3.415 5.12 4.84 ;
      RECT 4.89 1.82 5.235 3.245 ;
      RECT 5.865 1.82 6.195 3.245 ;
      RECT 0 -0.085 7.2 0.085 ;
      RECT 6.765 0.085 7.075 1.13 ;
      RECT 3.115 0.085 3.445 1.13 ;
      RECT 3.975 0.085 4.305 1.05 ;
      RECT 4.91 0.085 5.24 1.13 ;
      RECT 2.02 0.085 2.35 1.13 ;
      RECT 5.865 0.085 6.195 1.13 ;
      RECT 3.68 3.185 3.85 4.235 ;
      RECT 3.615 1.22 4.665 1.39 ;
      RECT 3.615 0.35 3.805 1.22 ;
      RECT 4.475 0.35 4.665 1.22 ;
      RECT 4.39 4.405 4.72 4.84 ;
      RECT 3.68 4.235 4.72 4.405 ;
      RECT 4.39 3.695 4.72 4.235 ;
      RECT 4.02 1.39 4.19 3.015 ;
      RECT 3.68 3.015 4.19 3.185 ;
      RECT 3.145 5.19 5.19 5.36 ;
      RECT 4.6 5.01 5.19 5.19 ;
      RECT 4.005 5.36 4.195 6.31 ;
      RECT 3.145 5.36 3.335 6.31 ;
      RECT 5.205 5.53 5.55 6.31 ;
      RECT 5.36 3.915 5.55 5.53 ;
      RECT 5.36 3.585 6.41 3.915 ;
      RECT 3.06 4.77 3.73 5.02 ;
      RECT 3.06 2.98 3.3 4.77 ;
      RECT 2.56 2.74 3.3 2.98 ;
      RECT 2.56 0.735 2.8 2.74 ;
      RECT 0 3.245 1.89 3.415 ;
    LAYER mcon ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 6.395 6.575 6.565 6.745 ;
      RECT 6.875 6.575 7.045 6.745 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 0.155 6.575 0.325 6.745 ;
      RECT 0.635 6.575 0.805 6.745 ;
      RECT 1.115 6.575 1.285 6.745 ;
      RECT 1.595 6.575 1.765 6.745 ;
      RECT 1.42 2.725 1.59 2.895 ;
      RECT 1.78 2.725 1.95 2.895 ;
      RECT 2.075 6.575 2.245 6.745 ;
      RECT 2.555 6.575 2.725 6.745 ;
      RECT 3.035 6.575 3.205 6.745 ;
      RECT 3.515 6.575 3.685 6.745 ;
      RECT 3.995 6.575 4.165 6.745 ;
      RECT 4.475 6.575 4.645 6.745 ;
      RECT 4.955 6.575 5.125 6.745 ;
      RECT 5.435 6.575 5.605 6.745 ;
      RECT 5.915 6.575 6.085 6.745 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.14 2.715 2.31 2.885 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
  END
END scs8ls_lpflow_lsbuf_lh_isowell_4

MACRO scs8ls_lpflow_isobufsrckapwr_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 14.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.065 1.43 2.725 1.695 ;
        RECT 0.925 1.695 4.305 1.865 ;
        RECT 0.925 1.43 1.255 1.695 ;
        RECT 4.045 1.22 4.305 1.695 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END SLEEP

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.345 0.415 1.76 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.4 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.4 0.245 ;
    END
  END vgnd

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.23 1.92 13.81 2.15 ;
    END
    ANTENNADIFFAREA 3.6288 ;
  END X

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 14.33 2.945 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.395 2.715 10.565 2.885 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.515 2.715 9.685 2.885 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.61 2.715 8.78 2.885 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.71 2.715 7.88 2.885 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.88 2.715 7.05 2.885 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.9 2.715 6.07 2.885 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 6.515 1.21 6.685 1.38 ;
      RECT 13.11 1.21 13.28 1.38 ;
      RECT 12.18 1.21 12.35 1.38 ;
      RECT 11.3 1.21 11.47 1.38 ;
      RECT 10.395 1.21 10.565 1.38 ;
      RECT 9.505 1.21 9.675 1.38 ;
      RECT 8.595 1.21 8.765 1.38 ;
      RECT 13.58 1.95 13.75 2.12 ;
      RECT 12.66 1.95 12.83 2.12 ;
      RECT 11.735 1.95 11.905 2.12 ;
      RECT 10.855 1.95 11.025 2.12 ;
      RECT 9.945 1.95 10.115 2.12 ;
      RECT 9.045 1.95 9.215 2.12 ;
      RECT 8.14 1.95 8.31 2.12 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.875 1.21 7.045 1.38 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.955 2.715 5.125 2.885 ;
      RECT 7.29 1.95 7.46 2.12 ;
      RECT 7.72 1.21 7.89 1.38 ;
      RECT 12.21 2.715 12.38 2.885 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 13.12 2.715 13.29 2.885 ;
      RECT 14.05 2.715 14.22 2.885 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.315 2.715 11.485 2.885 ;
    LAYER met1 ;
      RECT 6.455 1.18 13.34 1.41 ;
    LAYER li1 ;
      RECT 0.69 0.085 1.02 0.835 ;
      RECT 0 -0.085 14.4 0.085 ;
      RECT 1.63 0.085 1.96 0.58 ;
      RECT 2.49 0.085 2.82 0.58 ;
      RECT 3.35 0.085 3.68 0.58 ;
      RECT 4.23 0.085 4.56 0.58 ;
      RECT 4.915 0.085 5.165 0.81 ;
      RECT 5.775 0.085 6.025 0.81 ;
      RECT 6.655 0.085 6.985 0.81 ;
      RECT 7.655 0.085 7.865 0.745 ;
      RECT 8.5 0.085 8.735 0.745 ;
      RECT 9.415 0.085 9.68 0.745 ;
      RECT 10.33 0.085 10.605 0.745 ;
      RECT 11.235 0.085 11.515 0.745 ;
      RECT 12.11 0.085 12.445 0.745 ;
      RECT 13.05 0.085 13.355 0.745 ;
      RECT 13.965 0.085 14.285 0.745 ;
      RECT 1.075 2.575 1.325 3 ;
      RECT 1.075 2.405 3.215 2.575 ;
      RECT 2.145 2.575 2.315 2.995 ;
      RECT 3.045 2.575 3.215 2.75 ;
      RECT 3.045 2.375 3.215 2.405 ;
      RECT 1.075 2.035 1.335 2.405 ;
      RECT 3.045 2.75 4.125 2.92 ;
      RECT 3.935 2.375 4.125 2.75 ;
      RECT 0.585 1.175 3.635 1.26 ;
      RECT 3.305 1.26 3.635 1.515 ;
      RECT 0.26 1.09 3.635 1.175 ;
      RECT 0.1 2.1 0.37 3.075 ;
      RECT 0.1 1.93 0.755 2.1 ;
      RECT 0.585 1.26 0.755 1.93 ;
      RECT 0.26 1.005 0.785 1.09 ;
      RECT 0.26 0.255 0.52 1.005 ;
      RECT 1.565 1.26 1.895 1.515 ;
      RECT 6.8 2.29 7.05 2.98 ;
      RECT 5.37 2.12 5.7 2.98 ;
      RECT 5.37 1.95 6.655 2.12 ;
      RECT 6.27 2.12 6.6 2.98 ;
      RECT 6.485 1.46 6.655 1.95 ;
      RECT 6.485 1.15 7.09 1.46 ;
      RECT 5.345 1.13 7.09 1.15 ;
      RECT 5.345 0.98 6.935 1.13 ;
      RECT 5.345 0.395 5.595 0.98 ;
      RECT 6.225 0.395 6.475 0.98 ;
      RECT 13.97 1.82 14.28 2.98 ;
      RECT 7.665 1.19 7.945 1.52 ;
      RECT 8.515 1.19 8.835 1.52 ;
      RECT 9.435 1.19 9.74 1.52 ;
      RECT 10.325 1.19 10.63 1.52 ;
      RECT 11.23 1.19 11.53 1.52 ;
      RECT 12.11 1.19 12.43 1.52 ;
      RECT 13.05 1.19 13.345 1.52 ;
      RECT 11.705 0.395 11.93 2.98 ;
      RECT 11.245 1.82 11.515 2.98 ;
      RECT 10.82 0.745 11.05 2.98 ;
      RECT 10.775 0.395 11.05 0.745 ;
      RECT 10.345 1.82 10.64 2.98 ;
      RECT 9.92 0.745 10.145 2.98 ;
      RECT 9.85 0.395 10.145 0.745 ;
      RECT 9.43 1.82 9.725 2.98 ;
      RECT 9.015 0.745 9.245 2.98 ;
      RECT 8.915 0.395 9.245 0.745 ;
      RECT 8.53 1.82 8.83 2.98 ;
      RECT 8.125 0.745 8.33 2.98 ;
      RECT 8.045 0.395 8.33 0.745 ;
      RECT 7.665 1.82 7.935 2.98 ;
      RECT 13.525 0.395 13.775 2.98 ;
      RECT 13.05 1.82 13.345 2.98 ;
      RECT 12.63 0.395 12.87 2.98 ;
      RECT 12.13 1.82 12.45 2.98 ;
      RECT 5.9 2.29 6.07 2.98 ;
      RECT 4.92 1.95 5.17 2.98 ;
      RECT 7.26 0.745 7.485 2.98 ;
      RECT 7.2 0.395 7.485 0.745 ;
      RECT 1.615 2.035 4.7 2.205 ;
      RECT 4.475 1.78 4.7 2.035 ;
      RECT 4.475 1.35 6.315 1.78 ;
      RECT 4.475 0.92 4.7 1.35 ;
      RECT 1.2 0.75 4.7 0.92 ;
      RECT 1.615 2.205 1.945 2.235 ;
      RECT 1.2 0.645 1.46 0.75 ;
      RECT 3.415 2.205 3.745 2.58 ;
      RECT 2.13 0.645 2.32 0.75 ;
      RECT 2.99 0.625 3.18 0.75 ;
      RECT 3.86 0.625 4.03 0.75 ;
      RECT 0 3.245 14.4 3.415 ;
      RECT 2.515 2.745 2.845 3.245 ;
      RECT 4.315 2.375 4.645 3.245 ;
      RECT 0.555 2.27 0.835 3.245 ;
  END
END scs8ls_lpflow_isobufsrckapwr_16

MACRO scs8ls_lpflow_bleeder_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN short
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.25 1.78 2.175 ;
    END
    ANTENNAGATEAREA 0.315 ;
  END short

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.095 0.085 0.425 1.05 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 0 3.245 2.4 3.415 ;
      RECT 1.965 0.72 2.295 3.245 ;
    LAYER mcon ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_lpflow_bleeder_1

MACRO scs8ls_lpflow_fill_novpwr
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 0.48 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 0.48 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 0.48 0.085 ;
    LAYER mcon ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_lpflow_fill_novpwr

MACRO scs8ls_lpflow_sleep_aopwr_pargate
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.105 0.41 4.715 2.92 ;
    END
    ANTENNAGATEAREA 3.24 ;
  END sleep

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN aopwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 3.38 0 4.06 3.33 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.705 4.73 2.945 ;
        RECT 0.07 2.675 0.78 2.69 ;
        RECT 0.07 2.69 0.795 2.705 ;
        RECT 1.74 2.675 2.45 2.69 ;
        RECT 1.725 2.69 2.465 2.705 ;
        RECT 3.38 2.675 4.73 2.69 ;
        RECT 3.365 2.69 4.73 2.705 ;
    END
    PORT
      LAYER via ;
        RECT 3.855 0.44 4.005 0.59 ;
        RECT 3.855 2.74 4.005 2.89 ;
        RECT 3.435 0.44 3.585 0.59 ;
        RECT 3.435 2.74 3.585 2.89 ;
    END
  END aopwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 1.74 0 2.42 3.33 ;
    END
  END kapwr

  PIN realvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 2.56 0 3.24 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.92 0 1.6 3.33 ;
    END
    PORT
      LAYER via ;
        RECT 3.03 0.78 3.18 0.93 ;
        RECT 3.005 2.36 3.155 2.51 ;
        RECT 2.675 0.78 2.825 0.93 ;
        RECT 2.645 2.36 2.795 2.51 ;
        RECT 1.395 0.78 1.545 0.93 ;
        RECT 1.395 2.36 1.545 2.51 ;
        RECT 0.975 0.78 1.125 0.93 ;
        RECT 0.975 2.36 1.125 2.51 ;
    END
  END realvpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 0.89 0.785 3.265 0.985 ;
      RECT 2.59 0.725 3.265 0.755 ;
      RECT 2.56 0.755 3.265 0.785 ;
      RECT 0.89 0.71 1.63 0.745 ;
      RECT 0.89 0.745 1.665 0.78 ;
      RECT 0.89 0.78 1.7 0.785 ;
      RECT 3.405 0.665 4.09 0.675 ;
      RECT 1.77 0.385 4.09 0.585 ;
      RECT 3.365 0.585 4.09 0.625 ;
      RECT 3.405 0.625 4.09 0.665 ;
      RECT 1.77 0.585 2.5 0.615 ;
      RECT 1.77 0.615 2.47 0.645 ;
      RECT 0.89 2.305 3.27 2.535 ;
      RECT 0.89 2.535 1.66 2.55 ;
      RECT 0.89 2.55 1.645 2.565 ;
      RECT 2.545 2.535 3.27 2.55 ;
      RECT 2.56 2.55 3.27 2.565 ;
    LAYER li1 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 0.465 2.905 3.935 3.075 ;
      RECT 0.465 2.195 0.895 2.905 ;
      RECT 1.865 1.925 2.42 2.905 ;
      RECT 3.405 1.925 3.935 2.905 ;
      RECT 0.465 1.925 1.105 2.195 ;
      RECT 0.465 1.355 0.635 1.925 ;
      RECT 0.465 1.08 1.105 1.355 ;
      RECT 0.465 0.405 0.915 1.08 ;
      RECT 0.465 0.175 3.935 0.405 ;
      RECT 1.865 0.405 2.42 1.355 ;
      RECT 3.405 0.405 3.935 1.355 ;
      RECT 1.085 2.365 1.695 2.705 ;
      RECT 1.275 1.755 1.695 2.365 ;
      RECT 0.805 1.525 3.855 1.755 ;
      RECT 2.59 1.755 3.235 2.705 ;
      RECT 1.275 0.91 1.695 1.525 ;
      RECT 2.59 0.575 3.235 1.525 ;
      RECT 1.085 0.575 1.695 0.91 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.765 0.445 3.935 0.615 ;
      RECT 3.765 2.715 3.935 2.885 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.405 0.445 3.575 0.615 ;
      RECT 3.405 2.715 3.575 2.885 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.035 0.77 3.205 0.94 ;
      RECT 3.04 2.35 3.21 2.52 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.65 0.77 2.82 0.94 ;
      RECT 2.59 2.35 2.76 2.52 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.225 0.445 2.395 0.615 ;
      RECT 2.225 2.715 2.395 2.885 ;
      RECT 1.865 0.445 2.035 0.615 ;
      RECT 1.865 2.715 2.035 2.885 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.445 0.785 1.615 0.955 ;
      RECT 1.445 2.365 1.615 2.535 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.085 0.74 1.255 0.91 ;
      RECT 1.085 2.365 1.255 2.535 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_sleep_aopwr_pargate

MACRO scs8ls_lpflow_sleep_aopwr_pargate_2
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.105 0.41 8.53 2.92 ;
    END
    ANTENNAGATEAREA 7.56 ;
  END sleep

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN aopwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 3.555 0 4.325 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 7.195 0 7.965 3.33 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 8.57 2.945 ;
        RECT 1.705 2.655 2.535 2.675 ;
        RECT 3.525 2.655 4.355 2.675 ;
        RECT 5.345 2.655 6.175 2.675 ;
        RECT 7.165 2.655 7.995 2.675 ;
    END
    PORT
      LAYER via ;
        RECT 3.61 2.71 3.76 2.86 ;
        RECT 4.12 2.71 4.27 2.86 ;
        RECT 7.25 2.71 7.4 2.86 ;
        RECT 7.76 2.71 7.91 2.86 ;
        RECT 7.73 0.44 7.88 0.59 ;
        RECT 7.28 0.44 7.43 0.59 ;
        RECT 4.09 0.44 4.24 0.59 ;
        RECT 3.64 0.44 3.79 0.59 ;
    END
  END aopwr

  PIN realvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 0.805 0 1.595 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 6.285 0 7.055 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.465 0 5.235 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 2.645 0 3.415 3.33 ;
    END
    PORT
      LAYER via ;
        RECT 6.34 2.33 6.49 2.48 ;
        RECT 6.85 2.33 7 2.48 ;
        RECT 4.52 2.33 4.67 2.48 ;
        RECT 4.55 0.78 4.7 0.93 ;
        RECT 5.03 2.33 5.18 2.48 ;
        RECT 5 0.78 5.15 0.93 ;
        RECT 6.37 0.78 6.52 0.93 ;
        RECT 6.82 0.78 6.97 0.93 ;
        RECT 3.18 0.78 3.33 0.93 ;
        RECT 3.21 2.33 3.36 2.48 ;
        RECT 2.73 0.78 2.88 0.93 ;
        RECT 2.7 2.33 2.85 2.48 ;
        RECT 1.36 0.78 1.51 0.93 ;
        RECT 1.39 2.33 1.54 2.48 ;
        RECT 0.86 0.78 1.01 0.93 ;
        RECT 0.86 2.33 1.01 2.48 ;
    END
  END realvpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 1.735 0 2.505 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 5.375 0 6.145 3.33 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 1.735 0.585 2.505 0.645 ;
      RECT 1.735 0.385 7.965 0.585 ;
      RECT 3.555 0.585 4.325 0.645 ;
      RECT 5.375 0.585 6.145 0.645 ;
      RECT 7.195 0.585 7.965 0.645 ;
      RECT 0.775 2.515 1.625 2.535 ;
      RECT 0.775 2.245 7.085 2.515 ;
      RECT 2.615 2.515 3.445 2.535 ;
      RECT 4.435 2.515 5.265 2.535 ;
      RECT 6.255 2.515 7.085 2.535 ;
      RECT 0.775 0.785 7.055 0.985 ;
      RECT 0.775 0.725 1.595 0.785 ;
      RECT 2.645 0.725 3.415 0.785 ;
      RECT 4.465 0.725 5.235 0.785 ;
      RECT 6.285 0.725 7.055 0.785 ;
    LAYER li1 ;
      RECT 0.775 2.875 7.935 3.075 ;
      RECT 1.75 1.925 2.495 2.875 ;
      RECT 3.57 1.925 4.305 2.875 ;
      RECT 5.385 1.925 6.13 2.875 ;
      RECT 7.185 1.925 7.935 2.875 ;
      RECT 1.75 0.405 2.495 1.355 ;
      RECT 0.775 0.175 7.935 0.405 ;
      RECT 3.57 0.405 4.305 1.355 ;
      RECT 5.385 0.405 6.13 1.355 ;
      RECT 7.185 0.405 7.935 1.355 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 0.945 1.755 1.58 2.705 ;
      RECT 0.775 1.525 7.855 1.755 ;
      RECT 2.665 1.755 3.4 2.705 ;
      RECT 4.475 1.755 5.215 2.705 ;
      RECT 6.3 1.755 7.015 2.705 ;
      RECT 0.945 0.575 1.58 1.525 ;
      RECT 2.665 0.575 3.4 1.525 ;
      RECT 4.475 0.575 5.215 1.525 ;
      RECT 6.3 0.575 7.015 1.525 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 7.255 0.43 7.425 0.6 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.735 0.43 7.905 0.6 ;
      RECT 5.435 0.43 5.605 0.6 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 5.005 0.77 5.175 0.94 ;
      RECT 5.015 2.32 5.185 2.49 ;
      RECT 4.525 0.77 4.695 0.94 ;
      RECT 4.505 2.32 4.675 2.49 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 4.095 0.43 4.265 0.6 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.615 0.43 3.785 0.6 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 3.185 0.77 3.355 0.94 ;
      RECT 3.2 2.32 3.37 2.49 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 6.33 2.32 6.5 2.49 ;
      RECT 6.815 2.32 6.985 2.49 ;
      RECT 2.705 0.77 2.875 0.94 ;
      RECT 2.695 2.32 2.865 2.49 ;
      RECT 2.215 0.43 2.385 0.6 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.825 0.43 1.995 0.6 ;
      RECT 4.115 2.715 4.285 2.885 ;
      RECT 3.6 2.715 3.77 2.885 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.365 0.77 1.535 0.94 ;
      RECT 1.38 2.32 1.55 2.49 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.975 0.77 1.145 0.94 ;
      RECT 0.945 2.32 1.115 2.49 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 1.78 2.715 1.95 2.885 ;
      RECT 2.295 2.715 2.465 2.885 ;
      RECT 5.42 2.715 5.59 2.885 ;
      RECT 6.345 0.77 6.515 0.94 ;
      RECT 5.935 2.715 6.105 2.885 ;
      RECT 7.24 2.715 7.41 2.885 ;
      RECT 7.755 2.715 7.925 2.885 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 5.915 0.43 6.085 0.6 ;
      RECT 6.825 0.77 6.995 0.94 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
  END
END scs8ls_lpflow_sleep_aopwr_pargate_2

MACRO scs8ls_lpflow_sleep_aopwr_pargate_s8d
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.105 0.41 8.53 2.92 ;
    END
    ANTENNAGATEAREA 7.56 ;
  END sleep

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN realvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 5.3 0 6.88 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.75 0 3.33 3.33 ;
    END
    PORT
      LAYER via ;
        RECT 3.095 0.78 3.245 0.93 ;
        RECT 3.095 2.31 3.245 2.46 ;
        RECT 5.385 2.31 5.535 2.46 ;
        RECT 2.675 0.78 2.825 0.93 ;
        RECT 2.255 0.78 2.405 0.93 ;
        RECT 1.835 0.78 1.985 0.93 ;
        RECT 6.645 0.78 6.795 0.93 ;
        RECT 6.225 0.78 6.375 0.93 ;
        RECT 5.805 0.78 5.955 0.93 ;
        RECT 2.675 2.31 2.825 2.46 ;
        RECT 2.255 2.31 2.405 2.46 ;
        RECT 1.835 2.31 1.985 2.46 ;
        RECT 5.805 2.31 5.955 2.46 ;
        RECT 6.225 2.31 6.375 2.46 ;
        RECT 5.385 0.78 5.535 0.93 ;
        RECT 6.645 2.31 6.795 2.46 ;
    END
  END realvpwr

  PIN aopwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 7.02 0 8.035 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.47 0 4.245 3.33 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 8.57 2.945 ;
    END
    PORT
      LAYER via ;
        RECT 7.105 2.735 7.255 2.885 ;
        RECT 4.01 0.44 4.16 0.59 ;
        RECT 3.555 2.735 3.705 2.885 ;
        RECT 4.01 2.735 4.16 2.885 ;
        RECT 3.555 0.44 3.705 0.59 ;
        RECT 7.44 2.735 7.59 2.885 ;
        RECT 7.775 0.44 7.925 0.59 ;
        RECT 7.44 0.44 7.59 0.59 ;
        RECT 7.105 0.44 7.255 0.59 ;
        RECT 7.775 2.735 7.925 2.885 ;
    END
  END aopwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 0.62 0 1.61 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.385 0 5.16 3.33 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 1.75 2.255 6.88 2.515 ;
      RECT 0.6 0.585 1.61 0.645 ;
      RECT 0.6 0.385 8.035 0.585 ;
      RECT 3.47 0.585 5.16 0.645 ;
      RECT 7.02 0.585 8.035 0.645 ;
      RECT 1.75 0.785 6.88 0.985 ;
      RECT 1.75 0.725 3.33 0.785 ;
      RECT 5.3 0.725 6.88 0.785 ;
    LAYER li1 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 0.62 0.405 1.58 1.355 ;
      RECT 0.62 0.175 7.855 0.405 ;
      RECT 3.49 0.405 5.14 1.355 ;
      RECT 7.08 0.405 7.855 1.355 ;
      RECT 0.62 2.9 7.855 3.075 ;
      RECT 0.62 1.925 1.59 2.9 ;
      RECT 3.49 1.925 5.14 2.9 ;
      RECT 7.08 1.925 7.855 2.9 ;
      RECT 1.76 1.755 3.305 2.73 ;
      RECT 0.775 1.525 7.855 1.755 ;
      RECT 5.325 1.755 6.88 2.73 ;
      RECT 1.76 0.575 3.305 1.525 ;
      RECT 5.325 0.575 6.88 1.525 ;
    LAYER mcon ;
      RECT 6.215 2.3 6.385 2.47 ;
      RECT 1.81 2.3 1.98 2.47 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.38 0.43 1.55 0.6 ;
      RECT 1.02 0.43 1.19 0.6 ;
      RECT 2.245 2.3 2.415 2.47 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.66 0.43 0.83 0.6 ;
      RECT 2.665 2.3 2.835 2.47 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 6.65 2.3 6.82 2.47 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.215 0.77 6.385 0.94 ;
      RECT 0.66 2.725 0.83 2.895 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 6.65 0.77 6.82 0.94 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 5.795 0.77 5.965 0.94 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 7.66 0.43 7.83 0.6 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 4.93 0.43 5.1 0.6 ;
      RECT 5.36 0.77 5.53 0.94 ;
      RECT 1.38 2.725 1.55 2.895 ;
      RECT 4.93 2.725 5.1 2.895 ;
      RECT 4.46 2.725 4.63 2.895 ;
      RECT 4 2.725 4.17 2.895 ;
      RECT 3.53 2.725 3.7 2.895 ;
      RECT 1.02 2.725 1.19 2.895 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 7.66 2.725 7.83 2.895 ;
      RECT 7.1 2.725 7.27 2.895 ;
      RECT 4.46 0.43 4.63 0.6 ;
      RECT 4 0.43 4.17 0.6 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.53 0.43 3.7 0.6 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.1 0.77 3.27 0.94 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 2.665 0.77 2.835 0.94 ;
      RECT 3.1 2.3 3.27 2.47 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 5.36 2.3 5.53 2.47 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 2.245 0.77 2.415 0.94 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.81 0.77 1.98 0.94 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.795 2.3 5.965 2.47 ;
      RECT 7.1 0.43 7.27 0.6 ;
  END
END scs8ls_lpflow_sleep_aopwr_pargate_s8d

MACRO scs8ls_lpflow_sleep_kapwr_pargate_2
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.105 0.41 8.53 2.92 ;
    END
    ANTENNAGATEAREA 7.56 ;
  END sleep

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN aopwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 3.555 0 4.325 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 7.195 0 7.965 3.33 ;
    END
  END aopwr

  PIN realvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 0.805 0 1.595 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 6.285 0 7.055 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.465 0 5.235 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 2.645 0 3.415 3.33 ;
    END
    PORT
      LAYER via ;
        RECT 6.34 2.33 6.49 2.48 ;
        RECT 6.85 2.33 7 2.48 ;
        RECT 4.52 2.33 4.67 2.48 ;
        RECT 4.55 0.78 4.7 0.93 ;
        RECT 5.03 2.33 5.18 2.48 ;
        RECT 5 0.78 5.15 0.93 ;
        RECT 6.37 0.78 6.52 0.93 ;
        RECT 6.82 0.78 6.97 0.93 ;
        RECT 3.18 0.78 3.33 0.93 ;
        RECT 3.21 2.33 3.36 2.48 ;
        RECT 2.73 0.78 2.88 0.93 ;
        RECT 2.7 2.33 2.85 2.48 ;
        RECT 1.36 0.78 1.51 0.93 ;
        RECT 1.39 2.33 1.54 2.48 ;
        RECT 0.86 0.78 1.01 0.93 ;
        RECT 0.86 2.33 1.01 2.48 ;
    END
  END realvpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 1.735 0 2.505 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 5.375 0 6.145 3.33 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 8.57 2.945 ;
        RECT 1.705 2.655 2.535 2.675 ;
        RECT 3.525 2.655 4.355 2.675 ;
        RECT 5.345 2.655 6.175 2.675 ;
        RECT 7.165 2.655 7.995 2.675 ;
    END
    PORT
      LAYER via ;
        RECT 1.79 2.71 1.94 2.86 ;
        RECT 2.3 2.71 2.45 2.86 ;
        RECT 5.43 2.71 5.58 2.86 ;
        RECT 5.94 2.71 6.09 2.86 ;
        RECT 5.91 0.44 6.06 0.59 ;
        RECT 5.46 0.44 5.61 0.59 ;
        RECT 2.27 0.44 2.42 0.59 ;
        RECT 1.82 0.44 1.97 0.59 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 1.735 0.585 2.505 0.645 ;
      RECT 1.735 0.385 7.965 0.585 ;
      RECT 3.555 0.585 4.325 0.645 ;
      RECT 5.375 0.585 6.145 0.645 ;
      RECT 7.195 0.585 7.965 0.645 ;
      RECT 0.775 2.515 1.625 2.535 ;
      RECT 0.775 2.245 7.085 2.515 ;
      RECT 2.615 2.515 3.445 2.535 ;
      RECT 4.435 2.515 5.265 2.535 ;
      RECT 6.255 2.515 7.085 2.535 ;
      RECT 0.775 0.785 7.055 0.985 ;
      RECT 0.775 0.725 1.595 0.785 ;
      RECT 2.645 0.725 3.415 0.785 ;
      RECT 4.465 0.725 5.235 0.785 ;
      RECT 6.285 0.725 7.055 0.785 ;
    LAYER li1 ;
      RECT 0.775 2.875 7.935 3.075 ;
      RECT 1.75 1.925 2.495 2.875 ;
      RECT 3.57 1.925 4.305 2.875 ;
      RECT 5.385 1.925 6.13 2.875 ;
      RECT 7.185 1.925 7.935 2.875 ;
      RECT 1.75 0.405 2.495 1.355 ;
      RECT 0.775 0.175 7.935 0.405 ;
      RECT 3.57 0.405 4.305 1.355 ;
      RECT 5.385 0.405 6.13 1.355 ;
      RECT 7.185 0.405 7.935 1.355 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 0.945 1.755 1.58 2.705 ;
      RECT 0.775 1.525 7.855 1.755 ;
      RECT 2.665 1.755 3.4 2.705 ;
      RECT 4.475 1.755 5.215 2.705 ;
      RECT 6.3 1.755 7.015 2.705 ;
      RECT 0.945 0.575 1.58 1.525 ;
      RECT 2.665 0.575 3.4 1.525 ;
      RECT 4.475 0.575 5.215 1.525 ;
      RECT 6.3 0.575 7.015 1.525 ;
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 7.255 0.43 7.425 0.6 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.735 0.43 7.905 0.6 ;
      RECT 5.435 0.43 5.605 0.6 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 5.005 0.77 5.175 0.94 ;
      RECT 5.015 2.32 5.185 2.49 ;
      RECT 4.525 0.77 4.695 0.94 ;
      RECT 4.505 2.32 4.675 2.49 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 4.095 0.43 4.265 0.6 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.615 0.43 3.785 0.6 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 3.185 0.77 3.355 0.94 ;
      RECT 3.2 2.32 3.37 2.49 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 6.33 2.32 6.5 2.49 ;
      RECT 6.815 2.32 6.985 2.49 ;
      RECT 2.705 0.77 2.875 0.94 ;
      RECT 2.695 2.32 2.865 2.49 ;
      RECT 2.215 0.43 2.385 0.6 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.825 0.43 1.995 0.6 ;
      RECT 4.115 2.715 4.285 2.885 ;
      RECT 3.6 2.715 3.77 2.885 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.365 0.77 1.535 0.94 ;
      RECT 1.38 2.32 1.55 2.49 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.975 0.77 1.145 0.94 ;
      RECT 0.945 2.32 1.115 2.49 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 1.78 2.715 1.95 2.885 ;
      RECT 2.295 2.715 2.465 2.885 ;
      RECT 5.42 2.715 5.59 2.885 ;
      RECT 6.345 0.77 6.515 0.94 ;
      RECT 5.935 2.715 6.105 2.885 ;
      RECT 7.24 2.715 7.41 2.885 ;
      RECT 7.755 2.715 7.925 2.885 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 5.915 0.43 6.085 0.6 ;
      RECT 6.825 0.77 6.995 0.94 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
  END
END scs8ls_lpflow_sleep_kapwr_pargate_2

MACRO scs8ls_lpflow_sleep_kapwr_pargate_s8d
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.105 0.41 8.53 2.92 ;
    END
    ANTENNAGATEAREA 7.56 ;
  END sleep

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN realvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 5.3 0 6.88 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.75 0 3.33 3.33 ;
    END
    PORT
      LAYER via ;
        RECT 3.095 0.78 3.245 0.93 ;
        RECT 3.095 2.31 3.245 2.46 ;
        RECT 5.385 2.31 5.535 2.46 ;
        RECT 2.675 0.78 2.825 0.93 ;
        RECT 2.255 0.78 2.405 0.93 ;
        RECT 1.835 0.78 1.985 0.93 ;
        RECT 6.645 0.78 6.795 0.93 ;
        RECT 6.225 0.78 6.375 0.93 ;
        RECT 5.805 0.78 5.955 0.93 ;
        RECT 2.675 2.31 2.825 2.46 ;
        RECT 2.255 2.31 2.405 2.46 ;
        RECT 1.835 2.31 1.985 2.46 ;
        RECT 5.805 2.31 5.955 2.46 ;
        RECT 6.225 2.31 6.375 2.46 ;
        RECT 5.385 0.78 5.535 0.93 ;
        RECT 6.645 2.31 6.795 2.46 ;
    END
  END realvpwr

  PIN aopwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 7.02 0 8.035 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.47 0 4.245 3.33 ;
    END
  END aopwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 0.62 0 1.61 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.385 0 5.16 3.33 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 8.57 2.945 ;
    END
    PORT
      LAYER via ;
        RECT 0.705 2.735 0.855 2.885 ;
        RECT 4.925 0.44 5.075 0.59 ;
        RECT 4.925 2.735 5.075 2.885 ;
        RECT 4.47 2.735 4.62 2.885 ;
        RECT 4.47 0.44 4.62 0.59 ;
        RECT 1.04 2.735 1.19 2.885 ;
        RECT 1.375 0.44 1.525 0.59 ;
        RECT 1.04 0.44 1.19 0.59 ;
        RECT 0.705 0.44 0.855 0.59 ;
        RECT 1.375 2.735 1.525 2.885 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 1.75 2.255 6.88 2.515 ;
      RECT 0.6 0.585 1.61 0.645 ;
      RECT 0.6 0.385 8.035 0.585 ;
      RECT 3.47 0.585 5.16 0.645 ;
      RECT 7.02 0.585 8.035 0.645 ;
      RECT 1.75 0.785 6.88 0.985 ;
      RECT 1.75 0.725 3.33 0.785 ;
      RECT 5.3 0.725 6.88 0.785 ;
    LAYER li1 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 0.62 0.405 1.58 1.355 ;
      RECT 0.62 0.175 7.855 0.405 ;
      RECT 3.49 0.405 5.14 1.355 ;
      RECT 7.08 0.405 7.855 1.355 ;
      RECT 0.62 2.9 7.855 3.075 ;
      RECT 0.62 1.925 1.59 2.9 ;
      RECT 3.49 1.925 5.14 2.9 ;
      RECT 7.08 1.925 7.855 2.9 ;
      RECT 1.76 1.755 3.305 2.73 ;
      RECT 0.775 1.525 7.855 1.755 ;
      RECT 5.325 1.755 6.88 2.73 ;
      RECT 1.76 0.575 3.305 1.525 ;
      RECT 5.325 0.575 6.88 1.525 ;
    LAYER mcon ;
      RECT 6.215 2.3 6.385 2.47 ;
      RECT 1.81 2.3 1.98 2.47 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.38 0.43 1.55 0.6 ;
      RECT 1.02 0.43 1.19 0.6 ;
      RECT 2.245 2.3 2.415 2.47 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.66 0.43 0.83 0.6 ;
      RECT 2.665 2.3 2.835 2.47 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 6.65 2.3 6.82 2.47 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.215 0.77 6.385 0.94 ;
      RECT 0.66 2.725 0.83 2.895 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 6.65 0.77 6.82 0.94 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 5.795 0.77 5.965 0.94 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 7.66 0.43 7.83 0.6 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 4.93 0.43 5.1 0.6 ;
      RECT 5.36 0.77 5.53 0.94 ;
      RECT 1.38 2.725 1.55 2.895 ;
      RECT 4.93 2.725 5.1 2.895 ;
      RECT 4.46 2.725 4.63 2.895 ;
      RECT 4 2.725 4.17 2.895 ;
      RECT 3.53 2.725 3.7 2.895 ;
      RECT 1.02 2.725 1.19 2.895 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 7.66 2.725 7.83 2.895 ;
      RECT 7.1 2.725 7.27 2.895 ;
      RECT 4.46 0.43 4.63 0.6 ;
      RECT 4 0.43 4.17 0.6 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.53 0.43 3.7 0.6 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.1 0.77 3.27 0.94 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 2.665 0.77 2.835 0.94 ;
      RECT 3.1 2.3 3.27 2.47 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 5.36 2.3 5.53 2.47 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 2.245 0.77 2.415 0.94 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.81 0.77 1.98 0.94 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.795 2.3 5.965 2.47 ;
      RECT 7.1 0.43 7.27 0.6 ;
  END
END scs8ls_lpflow_sleep_kapwr_pargate_s8d

MACRO scs8ls_lpflow_sleep_pargate_s8d
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.105 0.41 8.53 2.92 ;
    END
    ANTENNAGATEAREA 7.56 ;
  END sleep

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN realvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 5.3 0 6.88 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.75 0 3.33 3.33 ;
    END
    PORT
      LAYER via ;
        RECT 3.095 0.78 3.245 0.93 ;
        RECT 3.095 2.33 3.245 2.48 ;
        RECT 5.385 2.33 5.535 2.48 ;
        RECT 2.675 0.78 2.825 0.93 ;
        RECT 2.255 0.78 2.405 0.93 ;
        RECT 1.835 0.78 1.985 0.93 ;
        RECT 6.645 0.78 6.795 0.93 ;
        RECT 6.225 0.78 6.375 0.93 ;
        RECT 5.805 0.78 5.955 0.93 ;
        RECT 2.675 2.33 2.825 2.48 ;
        RECT 2.255 2.33 2.405 2.48 ;
        RECT 1.835 2.33 1.985 2.48 ;
        RECT 5.805 2.33 5.955 2.48 ;
        RECT 6.225 2.33 6.375 2.48 ;
        RECT 5.385 0.78 5.535 0.93 ;
        RECT 6.645 2.33 6.795 2.48 ;
    END
  END realvpwr

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 7.02 0 8.035 3.49 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.47 0 4.245 3.49 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.385 0 5.16 3.49 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.62 0 1.61 3.49 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
    PORT
      LAYER via ;
        RECT 7.125 0.44 7.275 0.59 ;
        RECT 4.47 3.255 4.62 3.405 ;
        RECT 4.01 3.255 4.16 3.405 ;
        RECT 3.555 3.255 3.705 3.405 ;
        RECT 7.455 3.255 7.605 3.405 ;
        RECT 7.8 3.255 7.95 3.405 ;
        RECT 7.11 3.255 7.26 3.405 ;
        RECT 4.925 0.44 5.075 0.59 ;
        RECT 3.555 0.44 3.705 0.59 ;
        RECT 4.01 0.44 4.16 0.59 ;
        RECT 4.47 0.44 4.62 0.59 ;
        RECT 7.46 0.44 7.61 0.59 ;
        RECT 4.925 3.255 5.075 3.405 ;
        RECT 7.795 0.44 7.945 0.59 ;
        RECT 1.375 0.44 1.525 0.59 ;
        RECT 1.375 3.255 1.525 3.405 ;
        RECT 1.04 0.44 1.19 0.59 ;
        RECT 1.04 3.255 1.19 3.405 ;
        RECT 0.705 0.44 0.855 0.59 ;
        RECT 0.705 3.255 0.855 3.405 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 1.75 0.785 6.88 0.985 ;
      RECT 1.75 0.725 3.33 0.785 ;
      RECT 5.3 0.725 6.88 0.785 ;
      RECT 1.75 2.275 6.88 2.535 ;
      RECT 0.6 0.585 1.61 0.645 ;
      RECT 0.6 0.385 8.035 0.585 ;
      RECT 3.47 0.585 5.16 0.645 ;
      RECT 7.02 0.585 8.035 0.645 ;
    LAYER li1 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 0.795 2.9 7.855 3.245 ;
      RECT 0.795 1.95 1.59 2.9 ;
      RECT 3.49 1.95 5.14 2.9 ;
      RECT 7.08 1.95 7.855 2.9 ;
      RECT 0.62 0.43 1.58 1.38 ;
      RECT 0.62 0.2 7.855 0.43 ;
      RECT 3.49 0.43 5.14 1.38 ;
      RECT 7.08 0.43 7.855 1.38 ;
      RECT 1.76 1.78 3.305 2.73 ;
      RECT 0.775 1.55 7.855 1.78 ;
      RECT 5.325 1.78 6.88 2.73 ;
      RECT 1.76 0.6 3.305 1.55 ;
      RECT 5.325 0.6 6.88 1.55 ;
    LAYER mcon ;
      RECT 6.215 2.32 6.385 2.49 ;
      RECT 1.81 2.32 1.98 2.49 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.38 0.43 1.55 0.6 ;
      RECT 1.02 0.43 1.19 0.6 ;
      RECT 2.245 2.32 2.415 2.49 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.66 0.43 0.83 0.6 ;
      RECT 2.665 2.32 2.835 2.49 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 6.65 2.32 6.82 2.49 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.215 0.77 6.385 0.94 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 6.65 0.77 6.82 0.94 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 5.795 0.77 5.965 0.94 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 7.66 0.43 7.83 0.6 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 4.93 0.43 5.1 0.6 ;
      RECT 5.36 0.77 5.53 0.94 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 4.46 0.43 4.63 0.6 ;
      RECT 4 0.43 4.17 0.6 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.53 0.43 3.7 0.6 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.1 0.77 3.27 0.94 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 2.665 0.77 2.835 0.94 ;
      RECT 3.1 2.32 3.27 2.49 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 5.36 2.32 5.53 2.49 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 2.245 0.77 2.415 0.94 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.81 0.77 1.98 0.94 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.795 2.32 5.965 2.49 ;
      RECT 7.1 0.43 7.27 0.6 ;
  END
END scs8ls_lpflow_sleep_pargate_s8d

MACRO scs8ls_lpflow_sleep_vnwell_pargate
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.105 0.41 8.53 2.92 ;
    END
    ANTENNAGATEAREA 7.56 ;
  END sleep

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vnwell
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 8.57 2.945 ;
        RECT 1.705 2.655 2.535 2.675 ;
        RECT 3.525 2.655 4.355 2.675 ;
        RECT 5.345 2.655 6.175 2.675 ;
        RECT 7.165 2.655 7.995 2.675 ;
    END
  END vnwell

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN realvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 0.805 0 1.595 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 6.285 0 7.055 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.465 0 5.235 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 2.645 0 3.415 3.33 ;
    END
    PORT
      LAYER via ;
        RECT 6.34 2.33 6.49 2.48 ;
        RECT 6.85 2.33 7 2.48 ;
        RECT 4.52 2.33 4.67 2.48 ;
        RECT 4.55 0.78 4.7 0.93 ;
        RECT 5.03 2.33 5.18 2.48 ;
        RECT 5 0.78 5.15 0.93 ;
        RECT 6.37 0.78 6.52 0.93 ;
        RECT 6.82 0.78 6.97 0.93 ;
        RECT 3.18 0.78 3.33 0.93 ;
        RECT 3.21 2.33 3.36 2.48 ;
        RECT 2.73 0.78 2.88 0.93 ;
        RECT 2.7 2.33 2.85 2.48 ;
        RECT 1.36 0.78 1.51 0.93 ;
        RECT 1.39 2.33 1.54 2.48 ;
        RECT 0.86 0.78 1.01 0.93 ;
        RECT 0.86 2.33 1.01 2.48 ;
    END
  END realvpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 0.775 2.515 1.625 2.535 ;
      RECT 0.775 2.245 7.085 2.515 ;
      RECT 2.615 2.515 3.445 2.535 ;
      RECT 4.435 2.515 5.265 2.535 ;
      RECT 6.255 2.515 7.085 2.535 ;
      RECT 0.775 0.785 7.055 0.985 ;
      RECT 0.775 0.725 1.595 0.785 ;
      RECT 2.645 0.725 3.415 0.785 ;
      RECT 4.465 0.725 5.235 0.785 ;
      RECT 6.285 0.725 7.055 0.785 ;
      RECT 1.735 0.585 2.505 0.645 ;
      RECT 1.735 0.385 7.965 0.585 ;
      RECT 3.555 0.585 4.325 0.645 ;
      RECT 5.375 0.585 6.145 0.645 ;
      RECT 7.195 0.585 7.965 0.645 ;
    LAYER li1 ;
      RECT 2.665 0.575 3.4 2.705 ;
      RECT 0.775 2.875 7.935 3.075 ;
      RECT 1.75 0.405 2.495 2.875 ;
      RECT 3.57 0.405 4.305 2.875 ;
      RECT 5.385 0.405 6.13 2.875 ;
      RECT 7.185 0.405 7.935 2.875 ;
      RECT 0.775 0.175 7.935 0.405 ;
      RECT 0.825 0.575 1.58 2.705 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 6.3 0.575 7.015 2.705 ;
      RECT 4.475 0.575 5.215 2.705 ;
    LAYER mcon ;
      RECT 6.33 2.32 6.5 2.49 ;
      RECT 6.815 2.32 6.985 2.49 ;
      RECT 2.705 0.77 2.875 0.94 ;
      RECT 2.695 2.32 2.865 2.49 ;
      RECT 2.215 0.43 2.385 0.6 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.825 0.43 1.995 0.6 ;
      RECT 4.115 2.715 4.285 2.885 ;
      RECT 3.6 2.715 3.77 2.885 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.365 0.77 1.535 0.94 ;
      RECT 1.38 2.32 1.55 2.49 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.855 0.77 1.025 0.94 ;
      RECT 0.855 2.32 1.025 2.49 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 1.78 2.715 1.95 2.885 ;
      RECT 2.295 2.715 2.465 2.885 ;
      RECT 5.42 2.715 5.59 2.885 ;
      RECT 6.345 0.77 6.515 0.94 ;
      RECT 5.935 2.715 6.105 2.885 ;
      RECT 7.24 2.715 7.41 2.885 ;
      RECT 7.755 2.715 7.925 2.885 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 5.915 0.43 6.085 0.6 ;
      RECT 6.815 0.77 6.985 0.94 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 7.255 0.43 7.425 0.6 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.735 0.43 7.905 0.6 ;
      RECT 5.435 0.43 5.605 0.6 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 5.005 0.77 5.175 0.94 ;
      RECT 5.015 2.32 5.185 2.49 ;
      RECT 4.525 0.77 4.695 0.94 ;
      RECT 4.505 2.32 4.675 2.49 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 4.095 0.43 4.265 0.6 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.615 0.43 3.785 0.6 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 3.185 0.77 3.355 0.94 ;
      RECT 3.2 2.32 3.37 2.49 ;
      RECT 2.075 3.245 2.245 3.415 ;
  END
END scs8ls_lpflow_sleep_vnwell_pargate

MACRO scs8ls_lpflow_sleep_vnwell_pargate_s8d
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.105 0.41 8.53 2.92 ;
    END
    ANTENNAGATEAREA 7.56 ;
  END sleep

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vnwell
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 8.57 2.945 ;
    END
  END vnwell

  PIN realvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 5.3 0 6.88 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.75 0 3.33 3.33 ;
    END
    PORT
      LAYER via ;
        RECT 3.095 0.78 3.245 0.93 ;
        RECT 3.095 2.31 3.245 2.46 ;
        RECT 5.385 2.31 5.535 2.46 ;
        RECT 2.675 0.78 2.825 0.93 ;
        RECT 2.255 0.78 2.405 0.93 ;
        RECT 1.835 0.78 1.985 0.93 ;
        RECT 6.645 0.78 6.795 0.93 ;
        RECT 6.225 0.78 6.375 0.93 ;
        RECT 5.805 0.78 5.955 0.93 ;
        RECT 2.675 2.31 2.825 2.46 ;
        RECT 2.255 2.31 2.405 2.46 ;
        RECT 1.835 2.31 1.985 2.46 ;
        RECT 5.805 2.31 5.955 2.46 ;
        RECT 6.225 2.31 6.375 2.46 ;
        RECT 5.385 0.78 5.535 0.93 ;
        RECT 6.645 2.31 6.795 2.46 ;
    END
  END realvpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 1.75 2.255 6.88 2.515 ;
      RECT 0.6 0.585 1.61 0.645 ;
      RECT 0.6 0.385 8.035 0.585 ;
      RECT 3.47 0.585 5.16 0.645 ;
      RECT 7.02 0.585 8.035 0.645 ;
      RECT 1.75 0.785 6.88 0.985 ;
      RECT 1.75 0.725 3.33 0.785 ;
      RECT 5.3 0.725 6.88 0.785 ;
    LAYER li1 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 0.62 2.9 7.855 3.075 ;
      RECT 0.62 0.405 1.59 2.9 ;
      RECT 3.49 0.405 5.14 2.9 ;
      RECT 7.08 0.405 7.855 2.9 ;
      RECT 0.62 0.175 7.855 0.405 ;
      RECT 1.76 0.575 3.305 2.73 ;
      RECT 5.325 0.575 6.88 2.73 ;
    LAYER mcon ;
      RECT 6.215 0.77 6.385 0.94 ;
      RECT 0.66 2.725 0.83 2.895 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 6.65 0.77 6.82 0.94 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 5.795 0.77 5.965 0.94 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 7.66 0.43 7.83 0.6 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 4.93 0.43 5.1 0.6 ;
      RECT 5.36 0.77 5.53 0.94 ;
      RECT 1.38 2.725 1.55 2.895 ;
      RECT 4.93 2.725 5.1 2.895 ;
      RECT 4.46 2.725 4.63 2.895 ;
      RECT 4 2.725 4.17 2.895 ;
      RECT 3.53 2.725 3.7 2.895 ;
      RECT 1.02 2.725 1.19 2.895 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 7.66 2.725 7.83 2.895 ;
      RECT 7.1 2.725 7.27 2.895 ;
      RECT 4.46 0.43 4.63 0.6 ;
      RECT 4 0.43 4.17 0.6 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.53 0.43 3.7 0.6 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.1 0.77 3.27 0.94 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 2.665 0.77 2.835 0.94 ;
      RECT 3.1 2.3 3.27 2.47 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 5.36 2.3 5.53 2.47 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 2.245 0.77 2.415 0.94 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.81 0.77 1.98 0.94 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.795 2.3 5.965 2.47 ;
      RECT 7.1 0.43 7.27 0.6 ;
      RECT 6.215 2.3 6.385 2.47 ;
      RECT 1.81 2.3 1.98 2.47 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.38 0.43 1.55 0.6 ;
      RECT 1.02 0.43 1.19 0.6 ;
      RECT 2.245 2.3 2.415 2.47 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.66 0.43 0.83 0.6 ;
      RECT 2.665 2.3 2.835 2.47 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 6.65 2.3 6.82 2.47 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_sleep_vnwell_pargate_s8d

MACRO scs8ls_lpflow_sleep_fill_small
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 0.135 2.67 4.665 3.245 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_sleep_fill_small

MACRO scs8ls_lpflow_sleep_fill
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.135 2.67 8.505 3.245 ;
      RECT 0 3.245 8.64 3.415 ;
    LAYER mcon ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_sleep_fill

MACRO scs8ls_lpflow_isobufsrc_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 17.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.12 1.345 1.425 1.76 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END A

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2.295 1.55 16.67 1.78 ;
    END
    ANTENNAGATEAREA 4.464 ;
  END SLEEP

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2.975 1.92 15.875 2.15 ;
    END
    ANTENNADIFFAREA 6.3436 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 17.28 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 17.28 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 13.815 1.81 14.045 2.735 ;
      RECT 13.815 1.64 14.37 1.81 ;
      RECT 14.16 1.015 14.37 1.64 ;
      RECT 13.215 0.845 14.37 1.015 ;
      RECT 13.215 0.33 13.495 0.845 ;
      RECT 14.18 0.33 14.37 0.845 ;
      RECT 14.655 1.35 14.985 1.78 ;
      RECT 13.59 1.185 13.975 1.47 ;
      RECT 15.395 1.185 15.775 1.47 ;
      RECT 16.34 1.295 16.67 1.78 ;
      RECT 2.455 2.905 3.695 3.075 ;
      RECT 3.415 2.15 3.695 2.905 ;
      RECT 2.455 2.035 2.785 2.905 ;
      RECT 3.415 1.98 4.645 2.15 ;
      RECT 4.395 2.15 4.645 2.905 ;
      RECT 4.395 2.905 5.495 3.075 ;
      RECT 5.215 2.15 5.495 2.905 ;
      RECT 5.215 1.98 6.445 2.15 ;
      RECT 6.165 2.15 6.445 2.905 ;
      RECT 6.165 2.905 7.295 3.075 ;
      RECT 7.015 2.15 7.295 2.905 ;
      RECT 7.015 1.98 8.245 2.15 ;
      RECT 7.965 2.15 8.245 2.905 ;
      RECT 7.965 2.905 9.095 3.075 ;
      RECT 8.815 2.15 9.095 2.905 ;
      RECT 8.815 1.98 10.045 2.15 ;
      RECT 9.765 2.15 10.045 2.905 ;
      RECT 9.765 2.905 10.895 3.075 ;
      RECT 10.615 2.15 10.895 2.905 ;
      RECT 10.615 1.98 11.845 2.15 ;
      RECT 11.565 2.15 11.845 2.905 ;
      RECT 11.565 2.905 12.695 3.075 ;
      RECT 12.415 2.15 12.695 2.905 ;
      RECT 12.415 1.98 13.645 2.15 ;
      RECT 13.365 2.15 13.645 2.905 ;
      RECT 13.365 2.905 14.495 3.075 ;
      RECT 14.215 2.15 14.495 2.905 ;
      RECT 14.215 1.98 15.445 2.15 ;
      RECT 15.165 2.15 15.445 2.905 ;
      RECT 15.165 2.905 16.345 3.075 ;
      RECT 16.015 1.98 16.345 2.905 ;
      RECT 15.615 1.81 15.845 2.735 ;
      RECT 15.615 1.64 16.17 1.81 ;
      RECT 15.96 1.015 16.17 1.64 ;
      RECT 15.01 0.845 16.17 1.015 ;
      RECT 15.01 0.33 15.27 0.845 ;
      RECT 15.98 0.33 16.17 0.845 ;
      RECT 11.055 1.35 11.385 1.78 ;
      RECT 12.825 1.35 13.155 1.78 ;
      RECT 0.32 0.085 0.58 1.13 ;
      RECT 0 -0.085 17.28 0.085 ;
      RECT 1.18 0.085 1.44 0.835 ;
      RECT 2.04 0.085 2.37 0.835 ;
      RECT 2.98 0.085 3.31 0.675 ;
      RECT 3.84 0.085 4.1 1.125 ;
      RECT 4.7 0.085 5.03 0.675 ;
      RECT 5.59 0.085 5.845 1.125 ;
      RECT 6.48 0.085 6.81 0.675 ;
      RECT 7.34 0.085 7.625 1.125 ;
      RECT 8.28 0.085 8.61 0.675 ;
      RECT 9.16 0.085 9.425 1.125 ;
      RECT 10.08 0.085 10.41 0.675 ;
      RECT 10.945 0.085 11.23 1.125 ;
      RECT 11.88 0.085 12.21 0.675 ;
      RECT 12.76 0.085 13.035 1.125 ;
      RECT 13.68 0.085 14.01 0.675 ;
      RECT 14.54 0.085 14.83 1.125 ;
      RECT 15.48 0.085 15.81 0.675 ;
      RECT 16.34 0.085 16.67 1.125 ;
      RECT 0 3.245 17.28 3.415 ;
      RECT 3.865 2.32 4.195 3.245 ;
      RECT 5.665 2.32 5.995 3.245 ;
      RECT 7.465 2.32 7.795 3.245 ;
      RECT 9.265 2.32 9.595 3.245 ;
      RECT 11.065 2.32 11.395 3.245 ;
      RECT 12.865 2.32 13.195 3.245 ;
      RECT 14.665 2.32 14.995 3.245 ;
      RECT 1.005 2.27 1.335 3.245 ;
      RECT 1.935 2.27 2.265 3.245 ;
      RECT 16.515 1.95 16.795 3.245 ;
      RECT 0.105 1.93 0.38 3.245 ;
      RECT 5.625 1.35 5.955 1.78 ;
      RECT 10.215 1.81 10.445 2.735 ;
      RECT 10.215 1.64 10.775 1.81 ;
      RECT 10.56 1.015 10.775 1.64 ;
      RECT 9.615 0.845 10.775 1.015 ;
      RECT 9.615 0.33 9.895 0.845 ;
      RECT 10.58 0.33 10.775 0.845 ;
      RECT 12.015 1.81 12.245 2.735 ;
      RECT 12.015 1.64 12.57 1.81 ;
      RECT 12.36 1.015 12.57 1.64 ;
      RECT 11.41 0.845 12.57 1.015 ;
      RECT 11.41 0.33 11.67 0.845 ;
      RECT 12.38 0.33 12.57 0.845 ;
      RECT 4.815 1.81 5.045 2.735 ;
      RECT 4.815 1.64 5.405 1.81 ;
      RECT 5.17 1.015 5.405 1.64 ;
      RECT 4.27 0.845 5.405 1.015 ;
      RECT 4.27 0.33 4.53 0.845 ;
      RECT 5.21 0.33 5.405 0.845 ;
      RECT 10.025 1.185 10.375 1.47 ;
      RECT 11.8 1.185 12.165 1.47 ;
      RECT 4.655 1.185 4.985 1.47 ;
      RECT 9.21 1.35 9.575 1.78 ;
      RECT 6.445 1.185 6.775 1.47 ;
      RECT 7.455 1.35 7.785 1.78 ;
      RECT 6.615 1.81 6.845 2.735 ;
      RECT 6.615 1.64 7.17 1.81 ;
      RECT 6.96 1.015 7.17 1.64 ;
      RECT 6.015 0.845 7.17 1.015 ;
      RECT 6.015 0.33 6.295 0.845 ;
      RECT 6.98 0.33 7.17 0.845 ;
      RECT 3.895 1.35 4.225 1.78 ;
      RECT 2.965 1.81 3.245 2.735 ;
      RECT 2.965 1.64 3.67 1.81 ;
      RECT 3.45 1.015 3.67 1.64 ;
      RECT 2.55 0.845 3.67 1.015 ;
      RECT 2.55 0.33 2.81 0.845 ;
      RECT 3.48 0.33 3.67 0.845 ;
      RECT 8.415 1.81 8.645 2.735 ;
      RECT 8.415 1.64 8.97 1.81 ;
      RECT 8.76 1.015 8.97 1.64 ;
      RECT 7.81 0.845 8.97 1.015 ;
      RECT 7.81 0.33 8.07 0.845 ;
      RECT 8.78 0.33 8.97 0.845 ;
      RECT 2.925 1.185 3.255 1.47 ;
      RECT 2.295 1.35 2.605 1.865 ;
      RECT 8.22 1.185 8.58 1.47 ;
      RECT 0.59 2.1 0.835 2.98 ;
      RECT 0.59 1.93 2.125 2.1 ;
      RECT 1.505 2.1 1.765 2.98 ;
      RECT 1.595 1.175 2.125 1.93 ;
      RECT 0.75 1.005 2.125 1.175 ;
      RECT 0.75 0.35 1.01 1.005 ;
      RECT 1.61 0.35 1.87 1.005 ;
    LAYER mcon ;
      RECT 12.045 1.95 12.215 2.12 ;
      RECT 11.915 1.21 12.085 1.38 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 11.135 1.58 11.305 1.75 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.245 1.95 10.415 2.12 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.645 1.95 6.815 2.12 ;
      RECT 6.525 1.21 6.695 1.38 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.705 1.58 5.875 1.75 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.845 1.95 5.015 2.12 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 4.735 1.21 4.905 1.38 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 10.125 1.21 10.295 1.38 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.305 1.58 9.475 1.75 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 7.535 1.58 7.705 1.75 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.975 1.58 4.145 1.75 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.33 1.21 8.5 1.38 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 1.95 3.205 2.12 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.005 1.21 3.175 1.38 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.355 1.58 2.525 1.75 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.955 1.21 2.125 1.38 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 1.21 1.765 1.38 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.445 1.95 8.615 2.12 ;
      RECT 16.955 -0.085 17.125 0.085 ;
      RECT 16.955 3.245 17.125 3.415 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 16.44 1.58 16.61 1.75 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.645 1.95 15.815 2.12 ;
      RECT 15.525 1.21 15.695 1.38 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.735 1.58 14.905 1.75 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.845 1.95 14.015 2.12 ;
      RECT 13.725 1.21 13.895 1.38 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.905 1.58 13.075 1.75 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
    LAYER met1 ;
      RECT 1.535 1.18 15.755 1.41 ;
  END
END scs8ls_lpflow_isobufsrc_16

MACRO scs8ls_lpflow_isobufsrc_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.065 2.035 9.02 2.205 ;
        RECT 8.615 0.92 9.02 2.035 ;
        RECT 2.065 2.205 2.345 2.735 ;
        RECT 3.915 2.205 4.145 2.735 ;
        RECT 5.715 2.205 5.945 2.735 ;
        RECT 7.515 2.205 7.745 2.735 ;
        RECT 1.65 0.75 9.02 0.92 ;
        RECT 1.65 0.33 1.91 0.75 ;
        RECT 2.58 0.33 2.77 0.75 ;
        RECT 3.44 0.33 3.63 0.75 ;
        RECT 4.31 0.33 4.48 0.75 ;
        RECT 5.16 0.33 5.395 0.75 ;
        RECT 6.08 0.33 6.27 0.75 ;
        RECT 6.98 0.33 7.17 0.75 ;
        RECT 7.88 0.33 8.07 0.75 ;
    END
    ANTENNADIFFAREA 3.1052 ;
  END X

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.515 1.43 3.325 1.695 ;
        RECT 1.375 1.695 8.445 1.865 ;
        RECT 6.34 1.43 7.1 1.695 ;
        RECT 1.375 1.43 1.705 1.695 ;
        RECT 4.415 1.43 5.19 1.695 ;
        RECT 8.115 1.22 8.445 1.695 ;
    END
    ANTENNAGATEAREA 2.232 ;
  END SLEEP

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.345 0.865 1.76 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.12 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 9.12 0.085 ;
      RECT 8.24 0.085 8.91 0.58 ;
      RECT 0.28 0.085 0.54 1.13 ;
      RECT 1.14 0.085 1.47 0.835 ;
      RECT 2.08 0.085 2.41 0.58 ;
      RECT 2.94 0.085 3.27 0.58 ;
      RECT 3.8 0.085 4.13 0.58 ;
      RECT 4.66 0.085 4.99 0.58 ;
      RECT 5.58 0.085 5.91 0.58 ;
      RECT 6.44 0.085 6.77 0.58 ;
      RECT 7.38 0.085 7.71 0.58 ;
      RECT 0 3.245 9.12 3.415 ;
      RECT 8.415 2.375 8.99 3.245 ;
      RECT 1.035 2.27 1.365 3.245 ;
      RECT 0.105 1.93 0.38 3.245 ;
      RECT 2.965 2.715 3.295 3.245 ;
      RECT 4.765 2.715 5.095 3.245 ;
      RECT 6.565 2.715 6.895 3.245 ;
      RECT 7.065 2.905 8.245 3.075 ;
      RECT 7.915 2.375 8.245 2.905 ;
      RECT 1.555 2.035 1.885 2.905 ;
      RECT 1.555 2.905 2.795 3.075 ;
      RECT 2.515 2.545 2.795 2.905 ;
      RECT 2.515 2.375 3.745 2.545 ;
      RECT 3.495 2.545 3.745 2.905 ;
      RECT 3.495 2.905 4.595 3.075 ;
      RECT 4.315 2.545 4.595 2.905 ;
      RECT 4.315 2.375 5.545 2.545 ;
      RECT 5.265 2.545 5.545 2.905 ;
      RECT 5.265 2.905 6.395 3.075 ;
      RECT 6.115 2.545 6.395 2.905 ;
      RECT 6.115 2.375 7.345 2.545 ;
      RECT 7.065 2.545 7.345 2.905 ;
      RECT 1.035 1.175 7.77 1.26 ;
      RECT 7.44 1.26 7.77 1.525 ;
      RECT 0.71 1.09 7.77 1.175 ;
      RECT 0.55 2.1 0.865 2.98 ;
      RECT 0.55 1.93 1.205 2.1 ;
      RECT 1.035 1.26 1.205 1.93 ;
      RECT 0.71 1.005 1.235 1.09 ;
      RECT 0.71 0.35 0.97 1.005 ;
      RECT 2.015 1.26 2.345 1.515 ;
      RECT 3.755 1.26 4.085 1.515 ;
      RECT 5.595 1.26 5.925 1.525 ;
    LAYER mcon ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_isobufsrc_8

MACRO scs8ls_lpflow_sleep_kapwr_pargate
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.105 0.41 4.715 2.92 ;
    END
    ANTENNAGATEAREA 3.24 ;
  END sleep

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN aopwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 3.38 0 4.06 3.33 ;
    END
  END aopwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 1.74 0 2.42 3.33 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.705 4.73 2.945 ;
        RECT 0.07 2.675 0.78 2.69 ;
        RECT 0.07 2.69 0.795 2.705 ;
        RECT 1.74 2.675 2.45 2.69 ;
        RECT 1.725 2.69 2.465 2.705 ;
        RECT 3.38 2.675 4.73 2.69 ;
        RECT 3.365 2.69 4.73 2.705 ;
    END
    PORT
      LAYER via ;
        RECT 2.215 0.44 2.365 0.59 ;
        RECT 2.215 2.74 2.365 2.89 ;
        RECT 1.855 0.44 2.005 0.59 ;
        RECT 1.795 2.74 1.945 2.89 ;
    END
  END kapwr

  PIN realvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 2.56 0 3.24 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.92 0 1.6 3.33 ;
    END
    PORT
      LAYER via ;
        RECT 3.03 0.78 3.18 0.93 ;
        RECT 3.005 2.36 3.155 2.51 ;
        RECT 2.675 0.78 2.825 0.93 ;
        RECT 2.645 2.36 2.795 2.51 ;
        RECT 1.395 0.78 1.545 0.93 ;
        RECT 1.395 2.36 1.545 2.51 ;
        RECT 0.975 0.78 1.125 0.93 ;
        RECT 0.975 2.36 1.125 2.51 ;
    END
  END realvpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 0.89 0.785 3.265 0.985 ;
      RECT 2.59 0.725 3.265 0.755 ;
      RECT 2.56 0.755 3.265 0.785 ;
      RECT 0.89 0.71 1.63 0.745 ;
      RECT 0.89 0.745 1.665 0.78 ;
      RECT 0.89 0.78 1.7 0.785 ;
      RECT 3.405 0.665 4.09 0.675 ;
      RECT 1.77 0.385 4.09 0.585 ;
      RECT 3.365 0.585 4.09 0.625 ;
      RECT 3.405 0.625 4.09 0.665 ;
      RECT 1.77 0.585 2.5 0.615 ;
      RECT 1.77 0.615 2.47 0.645 ;
      RECT 0.89 2.305 3.27 2.535 ;
      RECT 0.89 2.535 1.66 2.55 ;
      RECT 0.89 2.55 1.645 2.565 ;
      RECT 2.545 2.535 3.27 2.55 ;
      RECT 2.56 2.55 3.27 2.565 ;
    LAYER li1 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 0.465 2.905 3.935 3.075 ;
      RECT 0.465 2.195 0.895 2.905 ;
      RECT 1.865 1.925 2.42 2.905 ;
      RECT 3.405 1.925 3.935 2.905 ;
      RECT 0.465 1.925 1.105 2.195 ;
      RECT 0.465 1.355 0.635 1.925 ;
      RECT 0.465 1.08 1.105 1.355 ;
      RECT 0.465 0.405 0.915 1.08 ;
      RECT 0.465 0.175 3.935 0.405 ;
      RECT 1.865 0.405 2.42 1.355 ;
      RECT 3.405 0.405 3.935 1.355 ;
      RECT 1.085 2.365 1.695 2.705 ;
      RECT 1.275 1.755 1.695 2.365 ;
      RECT 0.805 1.525 3.855 1.755 ;
      RECT 2.59 1.755 3.235 2.705 ;
      RECT 1.275 0.91 1.695 1.525 ;
      RECT 2.59 0.575 3.235 1.525 ;
      RECT 1.085 0.575 1.695 0.91 ;
    LAYER mcon ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.765 0.445 3.935 0.615 ;
      RECT 3.765 2.715 3.935 2.885 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.405 0.445 3.575 0.615 ;
      RECT 3.405 2.715 3.575 2.885 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.035 0.77 3.205 0.94 ;
      RECT 3.04 2.35 3.21 2.52 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.65 0.77 2.82 0.94 ;
      RECT 2.59 2.35 2.76 2.52 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.225 0.445 2.395 0.615 ;
      RECT 2.225 2.715 2.395 2.885 ;
      RECT 1.865 0.445 2.035 0.615 ;
      RECT 1.865 2.715 2.035 2.885 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.445 0.785 1.615 0.955 ;
      RECT 1.445 2.365 1.615 2.535 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.085 0.74 1.255 0.91 ;
      RECT 1.085 2.365 1.255 2.535 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_sleep_kapwr_pargate

MACRO scs8ls_lpflow_srsdfrtp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 21.12 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 20.205 0.35 20.525 1.99 ;
        RECT 20.205 1.99 20.505 2.98 ;
    END
    ANTENNADIFFAREA 0.5544 ;
  END Q

  PIN RESETB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.92 1.55 4.25 1.88 ;
    END
    ANTENNAGATEAREA 0.598 ;
  END RESETB

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.5 0.935 2.17 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.84 2.135 2.17 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.35 1.55 3.715 1.88 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 16.59 1.46 17.155 1.79 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END CLK

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.235 1.12 18.565 1.45 ;
    END
    ANTENNAGATEAREA 0.598 ;
  END SLEEPB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 21.12 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 21.12 3.575 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 21.05 2.945 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 20.315 -0.085 20.485 0.085 ;
      RECT 20.315 3.245 20.485 3.415 ;
      RECT 19.835 -0.085 20.005 0.085 ;
      RECT 20.795 3.245 20.965 3.415 ;
      RECT 20.795 -0.085 20.965 0.085 ;
      RECT 19.835 3.245 20.005 3.415 ;
      RECT 19.355 -0.085 19.525 0.085 ;
      RECT 19.355 3.245 19.525 3.415 ;
      RECT 18.875 -0.085 19.045 0.085 ;
      RECT 18.875 3.245 19.045 3.415 ;
      RECT 18.395 -0.085 18.565 0.085 ;
      RECT 18.395 3.245 18.565 3.415 ;
      RECT 17.915 -0.085 18.085 0.085 ;
      RECT 17.915 3.245 18.085 3.415 ;
      RECT 17.435 -0.085 17.605 0.085 ;
      RECT 17.435 2.735 17.605 2.905 ;
      RECT 17.435 3.245 17.605 3.415 ;
      RECT 16.955 -0.085 17.125 0.085 ;
      RECT 16.955 2.735 17.125 2.905 ;
      RECT 16.955 3.245 17.125 3.415 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 16.475 2.735 16.645 2.905 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 2.735 16.165 2.905 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 2.735 15.685 2.905 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 2.735 15.205 2.905 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 2.735 14.725 2.905 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
    LAYER li1 ;
      RECT 2.305 1.6 2.88 1.93 ;
      RECT 2.305 0.765 2.475 1.6 ;
      RECT 1.49 0.595 2.475 0.765 ;
      RECT 1.49 0.765 1.66 1.16 ;
      RECT 0.105 1.16 1.66 1.33 ;
      RECT 0.105 1.33 0.435 2.99 ;
      RECT 0.105 0.53 0.355 1.16 ;
      RECT 0 -0.085 21.12 0.085 ;
      RECT 20.695 0.085 20.965 1.13 ;
      RECT 18.805 0.085 19.055 0.805 ;
      RECT 19.855 0.085 20.025 1.13 ;
      RECT 0.535 0.085 0.865 0.99 ;
      RECT 3.615 0.085 3.865 1.04 ;
      RECT 7.05 0.085 7.38 0.835 ;
      RECT 8.02 0.085 8.35 0.825 ;
      RECT 11.365 0.085 11.695 0.985 ;
      RECT 13.125 0.085 13.455 0.81 ;
      RECT 17.475 0.085 17.805 0.61 ;
      RECT 0 3.245 21.12 3.415 ;
      RECT 20.695 1.82 20.965 3.245 ;
      RECT 6.12 2.77 6.45 3.245 ;
      RECT 7.85 2.605 8.18 3.245 ;
      RECT 3.245 2.41 4.3 3.245 ;
      RECT 19.715 1.815 20.035 3.245 ;
      RECT 0.645 2.34 0.975 3.245 ;
      RECT 18.735 1.815 18.985 2.18 ;
      RECT 18.735 1.145 18.905 1.815 ;
      RECT 18.735 0.975 19.685 1.145 ;
      RECT 19.515 1.145 19.685 1.315 ;
      RECT 19.235 0.345 19.685 0.975 ;
      RECT 19.515 1.315 19.94 1.645 ;
      RECT 12.21 2.35 19.325 2.52 ;
      RECT 19.155 1.645 19.325 2.35 ;
      RECT 19.075 1.315 19.345 1.645 ;
      RECT 9.835 2.565 12.54 2.735 ;
      RECT 12.21 2.52 12.54 2.565 ;
      RECT 9.835 2.04 10.5 2.565 ;
      RECT 10.19 0.605 10.5 2.04 ;
      RECT 13.625 2.52 13.955 2.97 ;
      RECT 16.25 1.74 16.42 2.35 ;
      RECT 15.985 1.41 16.42 1.74 ;
      RECT 17.895 1.85 18.49 2.18 ;
      RECT 16.93 0.78 18.345 0.95 ;
      RECT 18.015 0.345 18.345 0.78 ;
      RECT 17.895 0.95 18.065 1.85 ;
      RECT 16.93 0.425 17.1 0.78 ;
      RECT 14.985 0.255 17.1 0.425 ;
      RECT 14.985 0.425 15.315 0.6 ;
      RECT 14.015 0.6 15.315 0.77 ;
      RECT 14.015 0.77 14.185 1.32 ;
      RECT 12.93 1.32 14.185 1.5 ;
      RECT 14.525 2.69 17.73 3.025 ;
      RECT 16.855 2.01 17.495 2.18 ;
      RECT 17.325 1.29 17.495 2.01 ;
      RECT 16.59 1.12 17.495 1.29 ;
      RECT 16.105 1.11 16.76 1.12 ;
      RECT 14.355 0.95 16.76 1.11 ;
      RECT 14.355 1.11 14.525 1.67 ;
      RECT 14.355 0.94 16.435 0.95 ;
      RECT 11.64 1.67 14.525 1.84 ;
      RECT 16.105 0.595 16.435 0.94 ;
      RECT 11.64 1.51 11.97 1.67 ;
      RECT 11.1 2.01 16.08 2.18 ;
      RECT 14.695 1.93 16.08 2.01 ;
      RECT 11.1 1.325 11.43 2.01 ;
      RECT 14.695 1.28 14.955 1.93 ;
      RECT 11.1 1.155 12.235 1.325 ;
      RECT 11.905 0.575 12.235 1.155 ;
      RECT 12.695 0.98 13.845 1.15 ;
      RECT 12.695 0.575 12.945 0.98 ;
      RECT 13.675 0.575 13.845 0.98 ;
      RECT 8.555 2.905 13.455 3.075 ;
      RECT 8.555 2.825 8.725 2.905 ;
      RECT 13.125 2.745 13.455 2.905 ;
      RECT 8.395 2.435 8.725 2.825 ;
      RECT 5.78 2.43 8.725 2.435 ;
      RECT 5.78 2.435 7.68 2.6 ;
      RECT 7.51 2.265 8.725 2.43 ;
      RECT 4.925 2.6 5.95 2.77 ;
      RECT 8.395 1.665 8.725 2.265 ;
      RECT 4.925 1.92 5.095 2.6 ;
      RECT 8.395 1.495 9.4 1.665 ;
      RECT 4.885 1.59 5.215 1.92 ;
      RECT 9.07 1.665 9.4 1.825 ;
      RECT 8.395 1.335 8.99 1.495 ;
      RECT 7.32 1.845 8.135 2.095 ;
      RECT 7.965 1.175 8.135 1.845 ;
      RECT 6.28 1.165 8.135 1.175 ;
      RECT 6.28 1.175 6.61 1.485 ;
      RECT 6.28 1.005 9.53 1.165 ;
      RECT 9.2 1.165 9.53 1.285 ;
      RECT 7.59 0.995 9.53 1.005 ;
      RECT 7.59 0.575 7.84 0.995 ;
      RECT 9.2 0.435 9.53 0.995 ;
      RECT 9.2 0.265 10.93 0.435 ;
      RECT 10.68 0.435 10.93 2.395 ;
      RECT 5.265 2.26 5.555 2.43 ;
      RECT 5.265 2.09 7.11 2.26 ;
      RECT 6.78 1.675 7.11 2.09 ;
      RECT 5.385 1.265 5.555 2.09 ;
      RECT 6.78 1.345 7.795 1.675 ;
      RECT 5.375 0.935 5.555 1.265 ;
      RECT 4.615 0.425 4.865 1.08 ;
      RECT 4.615 0.255 6.59 0.425 ;
      RECT 6.26 0.425 6.59 0.835 ;
      RECT 2.305 2.1 4.755 2.24 ;
      RECT 4.47 2.24 4.755 2.99 ;
      RECT 2.98 2.07 4.715 2.1 ;
      RECT 4.545 1.42 4.715 2.07 ;
      RECT 4.545 1.25 5.205 1.42 ;
      RECT 5.035 0.765 5.205 1.25 ;
      RECT 5.035 0.595 6.055 0.765 ;
      RECT 5.725 0.765 6.055 1.265 ;
      RECT 1.96 2.51 2.635 2.99 ;
      RECT 1.225 2.34 2.635 2.51 ;
      RECT 2.305 2.325 2.635 2.34 ;
      RECT 2.305 2.24 3.08 2.325 ;
      RECT 1.225 1.5 2.08 1.67 ;
      RECT 1.83 0.935 2.08 1.5 ;
      RECT 1.225 1.67 1.395 2.34 ;
      RECT 2.645 1.21 4.375 1.38 ;
      RECT 2.645 0.74 2.975 1.21 ;
      RECT 4.045 0.58 4.375 1.21 ;
      RECT 1.07 0.425 1.32 0.99 ;
      RECT 1.07 0.255 3.405 0.425 ;
      RECT 3.155 0.425 3.405 1.04 ;
  END
END scs8ls_lpflow_srsdfrtp_2

MACRO scs8ls_lpflow_srsdfrtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 22.08 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 20.205 0.35 20.525 1.315 ;
        RECT 20.205 1.315 21.435 1.65 ;
        RECT 20.205 1.65 20.525 1.99 ;
        RECT 21.135 1.65 21.435 2.98 ;
        RECT 21.135 1.3 21.435 1.315 ;
        RECT 20.205 1.99 20.505 2.98 ;
        RECT 21.135 0.35 21.405 1.3 ;
    END
    ANTENNADIFFAREA 1.1532 ;
  END Q

  PIN RESETB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.92 1.55 4.25 1.88 ;
    END
    ANTENNAGATEAREA 0.598 ;
  END RESETB

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.5 0.935 2.17 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.84 2.135 2.17 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.35 1.55 3.715 1.88 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 16.59 1.46 17.155 1.79 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END CLK

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.235 1.12 18.565 1.45 ;
    END
    ANTENNAGATEAREA 0.598 ;
  END SLEEPB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 22.08 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 22.08 3.575 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 22.01 2.945 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.105 0.53 0.355 1.16 ;
      RECT 0 -0.085 22.08 0.085 ;
      RECT 21.575 0.085 21.855 1.13 ;
      RECT 18.805 0.085 19.075 0.805 ;
      RECT 19.855 0.085 20.025 1.13 ;
      RECT 20.695 0.085 20.965 1.13 ;
      RECT 0.535 0.085 0.865 0.99 ;
      RECT 3.615 0.085 3.865 1.04 ;
      RECT 7.05 0.085 7.38 0.835 ;
      RECT 8.02 0.085 8.35 0.825 ;
      RECT 11.365 0.085 11.695 0.985 ;
      RECT 13.125 0.085 13.455 0.81 ;
      RECT 17.475 0.085 17.805 0.61 ;
      RECT 0 3.245 22.08 3.415 ;
      RECT 21.605 1.82 21.885 3.245 ;
      RECT 6.12 2.77 6.45 3.245 ;
      RECT 7.85 2.605 8.18 3.245 ;
      RECT 3.245 2.41 4.3 3.245 ;
      RECT 19.715 1.815 20.035 3.245 ;
      RECT 20.695 1.82 20.965 3.245 ;
      RECT 0.645 2.34 0.975 3.245 ;
      RECT 18.735 1.815 18.985 2.18 ;
      RECT 18.735 1.145 18.905 1.815 ;
      RECT 18.735 0.975 19.685 1.145 ;
      RECT 19.515 1.145 19.685 1.315 ;
      RECT 19.245 0.345 19.685 0.975 ;
      RECT 19.515 1.315 19.94 1.645 ;
      RECT 12.21 2.35 19.325 2.52 ;
      RECT 19.155 1.645 19.325 2.35 ;
      RECT 19.075 1.315 19.345 1.645 ;
      RECT 9.835 2.565 12.54 2.735 ;
      RECT 12.21 2.52 12.54 2.565 ;
      RECT 9.835 2.04 10.5 2.565 ;
      RECT 10.19 0.605 10.5 2.04 ;
      RECT 13.625 2.52 13.955 2.97 ;
      RECT 16.25 1.74 16.42 2.35 ;
      RECT 15.985 1.41 16.42 1.74 ;
      RECT 17.895 1.85 18.49 2.18 ;
      RECT 16.93 0.78 18.345 0.95 ;
      RECT 18.015 0.345 18.345 0.78 ;
      RECT 17.895 0.95 18.065 1.85 ;
      RECT 16.93 0.425 17.1 0.78 ;
      RECT 14.985 0.255 17.1 0.425 ;
      RECT 14.985 0.425 15.315 0.6 ;
      RECT 14.015 0.6 15.315 0.77 ;
      RECT 14.015 0.77 14.185 1.32 ;
      RECT 12.93 1.32 14.185 1.5 ;
      RECT 14.525 2.69 17.73 3.025 ;
      RECT 16.855 2.01 17.495 2.18 ;
      RECT 17.325 1.29 17.495 2.01 ;
      RECT 16.59 1.12 17.495 1.29 ;
      RECT 16.105 1.11 16.76 1.12 ;
      RECT 14.355 0.95 16.76 1.11 ;
      RECT 14.355 1.11 14.525 1.67 ;
      RECT 14.355 0.94 16.435 0.95 ;
      RECT 11.64 1.67 14.525 1.84 ;
      RECT 16.105 0.595 16.435 0.94 ;
      RECT 11.64 1.51 11.97 1.67 ;
      RECT 11.1 2.01 16.08 2.18 ;
      RECT 14.695 1.93 16.08 2.01 ;
      RECT 11.1 1.325 11.43 2.01 ;
      RECT 14.695 1.28 14.955 1.93 ;
      RECT 11.1 1.155 12.235 1.325 ;
      RECT 11.905 0.575 12.235 1.155 ;
      RECT 12.695 0.98 13.845 1.15 ;
      RECT 12.695 0.575 12.945 0.98 ;
      RECT 13.675 0.575 13.845 0.98 ;
      RECT 8.555 2.905 13.455 3.075 ;
      RECT 8.555 2.825 8.725 2.905 ;
      RECT 13.125 2.745 13.455 2.905 ;
      RECT 8.395 2.435 8.725 2.825 ;
      RECT 5.78 2.43 8.725 2.435 ;
      RECT 5.78 2.435 7.68 2.6 ;
      RECT 7.51 2.265 8.725 2.43 ;
      RECT 4.925 2.6 5.95 2.77 ;
      RECT 8.395 1.665 8.725 2.265 ;
      RECT 4.925 1.92 5.095 2.6 ;
      RECT 8.395 1.495 9.4 1.665 ;
      RECT 4.885 1.59 5.215 1.92 ;
      RECT 9.07 1.665 9.4 1.825 ;
      RECT 8.395 1.335 8.99 1.495 ;
      RECT 7.32 1.845 8.135 2.095 ;
      RECT 7.965 1.175 8.135 1.845 ;
      RECT 6.28 1.165 8.135 1.175 ;
      RECT 6.28 1.175 6.61 1.485 ;
      RECT 6.28 1.005 9.53 1.165 ;
      RECT 9.2 1.165 9.53 1.285 ;
      RECT 7.59 0.995 9.53 1.005 ;
      RECT 7.59 0.575 7.84 0.995 ;
      RECT 9.2 0.435 9.53 0.995 ;
      RECT 9.2 0.265 10.93 0.435 ;
      RECT 10.68 0.435 10.93 2.395 ;
      RECT 5.265 2.26 5.555 2.43 ;
      RECT 5.265 2.09 7.11 2.26 ;
      RECT 6.78 1.675 7.11 2.09 ;
      RECT 5.385 1.265 5.555 2.09 ;
      RECT 6.78 1.345 7.795 1.675 ;
      RECT 5.375 0.935 5.555 1.265 ;
      RECT 4.615 0.425 4.865 1.08 ;
      RECT 4.615 0.255 6.59 0.425 ;
      RECT 6.26 0.425 6.59 0.835 ;
      RECT 2.305 2.1 4.755 2.24 ;
      RECT 4.47 2.24 4.755 2.99 ;
      RECT 2.98 2.07 4.715 2.1 ;
      RECT 4.545 1.42 4.715 2.07 ;
      RECT 4.545 1.25 5.205 1.42 ;
      RECT 5.035 0.765 5.205 1.25 ;
      RECT 5.035 0.595 6.055 0.765 ;
      RECT 5.725 0.765 6.055 1.265 ;
      RECT 1.96 2.51 2.635 2.99 ;
      RECT 1.225 2.34 2.635 2.51 ;
      RECT 2.305 2.325 2.635 2.34 ;
      RECT 2.305 2.24 3.08 2.325 ;
      RECT 1.225 1.5 2.08 1.67 ;
      RECT 1.83 0.935 2.08 1.5 ;
      RECT 1.225 1.67 1.395 2.34 ;
      RECT 2.645 1.21 4.375 1.38 ;
      RECT 2.645 0.74 2.975 1.21 ;
      RECT 4.045 0.58 4.375 1.21 ;
      RECT 1.07 0.425 1.32 0.99 ;
      RECT 1.07 0.255 3.405 0.425 ;
      RECT 3.155 0.425 3.405 1.04 ;
      RECT 2.305 1.6 2.88 1.93 ;
      RECT 2.305 0.765 2.475 1.6 ;
      RECT 1.49 0.595 2.475 0.765 ;
      RECT 1.49 0.765 1.66 1.16 ;
      RECT 0.105 1.16 1.66 1.33 ;
      RECT 0.105 1.33 0.435 2.99 ;
    LAYER mcon ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 16.955 -0.085 17.125 0.085 ;
      RECT 16.955 2.735 17.125 2.905 ;
      RECT 16.955 3.245 17.125 3.415 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 16.475 2.735 16.645 2.905 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 2.735 16.165 2.905 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 2.735 15.685 2.905 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 2.735 15.205 2.905 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 2.735 14.725 2.905 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 20.795 -0.085 20.965 0.085 ;
      RECT 20.795 3.245 20.965 3.415 ;
      RECT 20.315 -0.085 20.485 0.085 ;
      RECT 20.315 3.245 20.485 3.415 ;
      RECT 19.835 -0.085 20.005 0.085 ;
      RECT 21.275 3.245 21.445 3.415 ;
      RECT 21.275 -0.085 21.445 0.085 ;
      RECT 21.755 -0.085 21.925 0.085 ;
      RECT 21.755 3.245 21.925 3.415 ;
      RECT 19.835 3.245 20.005 3.415 ;
      RECT 19.355 -0.085 19.525 0.085 ;
      RECT 19.355 3.245 19.525 3.415 ;
      RECT 18.875 -0.085 19.045 0.085 ;
      RECT 18.875 3.245 19.045 3.415 ;
      RECT 18.395 -0.085 18.565 0.085 ;
      RECT 18.395 3.245 18.565 3.415 ;
      RECT 17.915 -0.085 18.085 0.085 ;
      RECT 17.915 3.245 18.085 3.415 ;
      RECT 17.435 -0.085 17.605 0.085 ;
      RECT 17.435 2.735 17.605 2.905 ;
      RECT 17.435 3.245 17.605 3.415 ;
  END
END scs8ls_lpflow_srsdfrtp_4

MACRO scs8ls_lpflow_srsdfstp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 19.2 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SETB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.725 0.78 7.16 1.03 ;
        RECT 6.725 1.03 7.22 1.265 ;
    END
    ANTENNAGATEAREA 0.439 ;
  END SETB

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.365 0.35 18.62 3.075 ;
    END
    ANTENNADIFFAREA 0.558 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.545 1.43 1.875 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.725 1.18 3.235 1.555 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.205 0.835 1.875 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.935 1.22 16.26 2.15 ;
    END
    ANTENNAGATEAREA 0.598 ;
  END SLEEPB

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 14.965 1.18 15.235 2.15 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END CLK

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 19.2 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 19.2 3.575 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 19.13 2.945 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 13.8 2.49 14.595 2.52 ;
      RECT 15.745 0.88 16.835 1.05 ;
      RECT 16.455 1.05 16.835 2.15 ;
      RECT 16.665 0.8 16.835 0.88 ;
      RECT 16.665 0.63 17.125 0.8 ;
      RECT 16.795 0.42 17.125 0.63 ;
      RECT 12.165 0.255 15.915 0.425 ;
      RECT 15.745 0.425 15.915 0.88 ;
      RECT 11.625 1.125 12.335 1.375 ;
      RECT 12.165 0.425 12.335 1.125 ;
      RECT 13.32 0.425 13.65 0.715 ;
      RECT 12.655 2.905 16.305 3.075 ;
      RECT 14.905 2.66 16.305 2.905 ;
      RECT 15.405 1.58 15.765 2.15 ;
      RECT 15.405 0.845 15.575 1.58 ;
      RECT 14.765 0.595 15.575 0.845 ;
      RECT 10.655 2.055 10.985 2.215 ;
      RECT 10.655 1.885 13.015 2.055 ;
      RECT 11.475 2.055 11.805 2.235 ;
      RECT 12.845 1.055 13.015 1.885 ;
      RECT 12.845 0.885 14.55 1.055 ;
      RECT 14.22 1.055 14.55 1.26 ;
      RECT 7.845 2.905 8.695 3.075 ;
      RECT 8.525 1.74 8.695 2.905 ;
      RECT 7.845 1.605 8.015 2.905 ;
      RECT 8.525 1.355 8.755 1.74 ;
      RECT 5.65 1.45 8.015 1.605 ;
      RECT 8.525 0.765 8.695 1.355 ;
      RECT 5.65 1.605 6.895 1.62 ;
      RECT 6.725 1.435 8.015 1.45 ;
      RECT 8.525 0.595 9.535 0.765 ;
      RECT 7.845 1.37 8.015 1.435 ;
      RECT 9.365 0.765 9.535 2.405 ;
      RECT 9.365 2.405 12.145 2.575 ;
      RECT 11.975 2.395 12.145 2.405 ;
      RECT 11.975 2.225 13.355 2.395 ;
      RECT 13.185 2.18 13.355 2.225 ;
      RECT 13.185 2.01 14.21 2.18 ;
      RECT 14.04 1.8 14.21 2.01 ;
      RECT 14.04 1.55 14.37 1.8 ;
      RECT 5.65 0.92 5.82 1.45 ;
      RECT 5.08 0.75 5.82 0.92 ;
      RECT 5.08 0.425 5.25 0.75 ;
      RECT 3.42 0.255 5.25 0.425 ;
      RECT 3.42 0.425 4.015 0.555 ;
      RECT 3.42 0.555 3.67 1.695 ;
      RECT 3.42 1.695 4.255 2.025 ;
      RECT 4.005 2.025 4.255 2.395 ;
      RECT 10.425 1.205 11.455 1.375 ;
      RECT 10.425 0.605 10.595 1.205 ;
      RECT 11.205 0.605 11.455 1.205 ;
      RECT 10.165 1.545 10.415 2.145 ;
      RECT 8.185 1.2 8.355 2.565 ;
      RECT 7.825 0.595 8.355 1.2 ;
      RECT 6.68 2.485 7.01 2.58 ;
      RECT 5.9 2.29 7.01 2.485 ;
      RECT 5.9 2.13 6.23 2.29 ;
      RECT 5.31 1.79 6.77 1.96 ;
      RECT 6.44 1.96 6.77 2.015 ;
      RECT 5.205 2.67 5.535 3 ;
      RECT 5.31 1.96 5.48 2.67 ;
      RECT 5.31 1.26 5.48 1.79 ;
      RECT 4.745 1.135 5.48 1.26 ;
      RECT 4.41 1.09 5.48 1.135 ;
      RECT 4.41 0.82 4.91 1.09 ;
      RECT 5.99 1.09 6.555 1.27 ;
      RECT 6.305 0.595 6.555 1.09 ;
      RECT 4.77 1.58 5.125 2.035 ;
      RECT 3.665 2.655 5.035 2.825 ;
      RECT 3.665 2.395 3.835 2.655 ;
      RECT 4.43 1.525 4.6 2.655 ;
      RECT 1.44 2.225 3.835 2.395 ;
      RECT 3.98 1.355 4.6 1.525 ;
      RECT 3.98 0.755 4.23 1.355 ;
      RECT 1.44 2.395 1.77 2.735 ;
      RECT 1.6 1.035 1.77 2.225 ;
      RECT 0.92 0.865 1.77 1.035 ;
      RECT 0.92 0.575 1.25 0.865 ;
      RECT 1.94 1.725 2.74 2.055 ;
      RECT 2.385 0.675 2.74 1.01 ;
      RECT 1.94 1.305 2.555 1.725 ;
      RECT 2.385 1.01 2.555 1.305 ;
      RECT 1.02 2.905 2.22 3.075 ;
      RECT 1.97 2.65 2.22 2.905 ;
      RECT 1.02 2.215 1.19 2.905 ;
      RECT 0.1 2.045 1.19 2.215 ;
      RECT 0.1 2.215 0.43 3.065 ;
      RECT 0 3.245 19.2 3.415 ;
      RECT 18.805 1.815 19.065 3.245 ;
      RECT 17.855 1.815 18.185 3.245 ;
      RECT 6.085 2.75 6.415 3.245 ;
      RECT 2.925 2.565 3.255 3.245 ;
      RECT 7.25 2.29 7.58 3.245 ;
      RECT 0.6 2.385 0.85 3.245 ;
      RECT 0 -0.085 19.2 0.085 ;
      RECT 18.79 0.085 19.05 1.015 ;
      RECT 7.33 0.085 7.5 0.895 ;
      RECT 10.775 0.085 11.025 1.035 ;
      RECT 11.745 0.085 11.995 0.955 ;
      RECT 16.085 0.085 16.335 0.71 ;
      RECT 17.86 0.085 18.19 1.015 ;
      RECT 0.1 0.085 0.43 1.035 ;
      RECT 1.94 0.085 2.19 1.035 ;
      RECT 2.92 0.085 3.25 1.01 ;
      RECT 5.465 0.085 5.795 0.58 ;
      RECT 17.39 1.995 17.675 2.675 ;
      RECT 17.505 1.55 17.675 1.995 ;
      RECT 17.505 1.22 18.18 1.55 ;
      RECT 17.505 0.675 17.675 1.22 ;
      RECT 17.325 0.35 17.675 0.675 ;
      RECT 13.8 2.35 17.22 2.49 ;
      RECT 14.425 2.32 17.22 2.35 ;
      RECT 17.05 1.825 17.22 2.32 ;
      RECT 17.005 1.495 17.335 1.825 ;
      RECT 8.925 2.745 12.485 3.075 ;
      RECT 12.315 2.735 12.485 2.745 ;
      RECT 8.925 2.235 9.195 2.745 ;
      RECT 12.315 2.565 14.13 2.735 ;
      RECT 8.925 1.225 9.095 2.235 ;
      RECT 13.8 2.52 14.13 2.565 ;
      RECT 8.865 0.935 9.195 1.225 ;
    LAYER mcon ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 2.735 16.165 2.905 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 1.58 15.685 1.75 ;
      RECT 15.515 2.735 15.685 2.905 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 2.735 15.205 2.905 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.24 1.58 10.41 1.75 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 1.58 5.125 1.75 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 18.395 -0.085 18.565 0.085 ;
      RECT 18.395 3.245 18.565 3.415 ;
      RECT 17.915 -0.085 18.085 0.085 ;
      RECT 17.915 3.245 18.085 3.415 ;
      RECT 17.435 -0.085 17.605 0.085 ;
      RECT 17.435 3.245 17.605 3.415 ;
      RECT 16.955 -0.085 17.125 0.085 ;
      RECT 16.955 3.245 17.125 3.415 ;
      RECT 18.875 3.245 19.045 3.415 ;
      RECT 18.875 -0.085 19.045 0.085 ;
    LAYER met1 ;
      RECT 4.895 1.735 5.185 1.78 ;
      RECT 4.895 1.595 15.745 1.735 ;
      RECT 10.18 1.735 10.47 1.78 ;
      RECT 15.455 1.735 15.745 1.78 ;
      RECT 4.895 1.55 5.185 1.595 ;
      RECT 10.18 1.55 10.47 1.595 ;
      RECT 15.455 1.55 15.745 1.595 ;
  END
END scs8ls_lpflow_srsdfstp_2

MACRO scs8ls_lpflow_srsdfstp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 20.16 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SETB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.725 0.78 7.16 1.03 ;
        RECT 6.725 1.03 7.22 1.265 ;
    END
    ANTENNAGATEAREA 0.439 ;
  END SETB

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.365 1.77 18.62 3.075 ;
        RECT 18.365 1.695 19.49 1.77 ;
        RECT 18.425 1.545 19.49 1.695 ;
        RECT 19.26 1.77 19.49 3.075 ;
        RECT 18.425 1.065 18.62 1.545 ;
        RECT 19.22 0.35 19.49 1.545 ;
        RECT 18.365 0.35 18.62 1.065 ;
    END
    ANTENNADIFFAREA 1.1531 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.545 1.43 1.875 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.725 1.18 3.235 1.555 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.205 0.835 1.875 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.935 1.22 16.26 2.15 ;
    END
    ANTENNAGATEAREA 0.598 ;
  END SLEEPB

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 14.965 1.18 15.235 2.15 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END CLK

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 20.16 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 20.16 3.575 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 20.09 2.945 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 12.845 1.055 13.015 1.885 ;
      RECT 12.845 0.885 14.55 1.055 ;
      RECT 14.22 1.055 14.55 1.26 ;
      RECT 7.845 2.905 8.695 3.075 ;
      RECT 8.525 1.74 8.695 2.905 ;
      RECT 7.845 1.605 8.015 2.905 ;
      RECT 8.525 1.355 8.755 1.74 ;
      RECT 5.65 1.45 8.015 1.605 ;
      RECT 8.525 0.765 8.695 1.355 ;
      RECT 5.65 1.605 6.895 1.62 ;
      RECT 6.725 1.435 8.015 1.45 ;
      RECT 8.525 0.595 9.535 0.765 ;
      RECT 7.845 1.37 8.015 1.435 ;
      RECT 9.365 0.765 9.535 2.405 ;
      RECT 9.365 2.405 12.145 2.575 ;
      RECT 11.975 2.395 12.145 2.405 ;
      RECT 11.975 2.225 13.355 2.395 ;
      RECT 13.185 2.18 13.355 2.225 ;
      RECT 13.185 2.01 14.21 2.18 ;
      RECT 14.04 1.8 14.21 2.01 ;
      RECT 14.04 1.55 14.37 1.8 ;
      RECT 5.65 0.92 5.82 1.45 ;
      RECT 5.08 0.75 5.82 0.92 ;
      RECT 5.08 0.425 5.25 0.75 ;
      RECT 3.42 0.255 5.25 0.425 ;
      RECT 3.42 0.425 4.015 0.555 ;
      RECT 3.42 0.555 3.67 1.695 ;
      RECT 3.42 1.695 4.255 2.025 ;
      RECT 4.005 2.025 4.255 2.395 ;
      RECT 10.425 1.205 11.455 1.375 ;
      RECT 10.425 0.605 10.595 1.205 ;
      RECT 11.205 0.605 11.455 1.205 ;
      RECT 10.165 1.545 10.415 2.145 ;
      RECT 8.185 1.2 8.355 2.565 ;
      RECT 7.825 0.595 8.355 1.2 ;
      RECT 6.68 2.485 7.01 2.58 ;
      RECT 5.9 2.29 7.01 2.485 ;
      RECT 5.9 2.13 6.23 2.29 ;
      RECT 5.31 1.79 6.77 1.96 ;
      RECT 6.44 1.96 6.77 2.015 ;
      RECT 5.205 2.67 5.535 3 ;
      RECT 5.31 1.96 5.48 2.67 ;
      RECT 5.31 1.26 5.48 1.79 ;
      RECT 4.745 1.135 5.48 1.26 ;
      RECT 4.41 1.09 5.48 1.135 ;
      RECT 4.41 0.82 4.91 1.09 ;
      RECT 5.99 1.09 6.555 1.27 ;
      RECT 6.305 0.595 6.555 1.09 ;
      RECT 4.77 1.58 5.125 2.035 ;
      RECT 3.665 2.655 5.035 2.825 ;
      RECT 3.665 2.395 3.835 2.655 ;
      RECT 4.43 1.525 4.6 2.655 ;
      RECT 1.44 2.225 3.835 2.395 ;
      RECT 3.98 1.355 4.6 1.525 ;
      RECT 3.98 0.755 4.23 1.355 ;
      RECT 1.44 2.395 1.77 2.735 ;
      RECT 1.6 1.035 1.77 2.225 ;
      RECT 0.92 0.865 1.77 1.035 ;
      RECT 0.92 0.575 1.25 0.865 ;
      RECT 1.94 1.725 2.74 2.055 ;
      RECT 2.385 0.675 2.74 1.01 ;
      RECT 1.94 1.305 2.555 1.725 ;
      RECT 2.385 1.01 2.555 1.305 ;
      RECT 1.02 2.905 2.22 3.075 ;
      RECT 1.97 2.65 2.22 2.905 ;
      RECT 1.02 2.215 1.19 2.905 ;
      RECT 0.1 2.045 1.19 2.215 ;
      RECT 0.1 2.215 0.43 3.065 ;
      RECT 0 -0.085 20.16 0.085 ;
      RECT 19.66 0.085 19.985 1.015 ;
      RECT 7.33 0.085 7.5 0.895 ;
      RECT 10.775 0.085 11.025 1.035 ;
      RECT 11.745 0.085 11.995 0.955 ;
      RECT 16.085 0.085 16.335 0.71 ;
      RECT 17.86 0.085 18.19 1.015 ;
      RECT 18.79 0.085 19.05 1 ;
      RECT 0.1 0.085 0.43 1.035 ;
      RECT 1.94 0.085 2.19 1.035 ;
      RECT 2.92 0.085 3.25 1.01 ;
      RECT 5.465 0.085 5.795 0.58 ;
      RECT 0 3.245 20.16 3.415 ;
      RECT 19.695 1.815 19.985 3.245 ;
      RECT 17.855 1.815 18.185 3.245 ;
      RECT 18.79 1.965 19.065 3.245 ;
      RECT 6.085 2.75 6.415 3.245 ;
      RECT 2.925 2.565 3.255 3.245 ;
      RECT 7.25 2.29 7.58 3.245 ;
      RECT 0.6 2.385 0.85 3.245 ;
      RECT 17.39 1.84 17.675 2.995 ;
      RECT 17.505 1.55 17.675 1.84 ;
      RECT 17.505 1.22 18.255 1.55 ;
      RECT 17.505 1.05 17.675 1.22 ;
      RECT 17.325 0.33 17.675 1.05 ;
      RECT 13.8 2.35 17.22 2.49 ;
      RECT 14.425 2.32 17.22 2.35 ;
      RECT 17.05 1.675 17.22 2.32 ;
      RECT 17.005 1.345 17.335 1.675 ;
      RECT 8.925 2.745 12.485 3.075 ;
      RECT 12.315 2.735 12.485 2.745 ;
      RECT 8.925 2.235 9.195 2.745 ;
      RECT 12.315 2.565 14.13 2.735 ;
      RECT 8.925 1.225 9.095 2.235 ;
      RECT 13.8 2.52 14.13 2.565 ;
      RECT 8.865 0.935 9.195 1.225 ;
      RECT 13.8 2.49 14.595 2.52 ;
      RECT 15.745 0.88 16.835 1.05 ;
      RECT 16.455 1.05 16.835 2.15 ;
      RECT 16.665 0.8 16.835 0.88 ;
      RECT 16.665 0.63 17.125 0.8 ;
      RECT 16.795 0.42 17.125 0.63 ;
      RECT 12.165 0.255 15.915 0.425 ;
      RECT 15.745 0.425 15.915 0.88 ;
      RECT 11.625 1.125 12.335 1.375 ;
      RECT 12.165 0.425 12.335 1.125 ;
      RECT 13.32 0.425 13.65 0.715 ;
      RECT 12.655 2.905 16.305 3.075 ;
      RECT 14.905 2.66 16.305 2.905 ;
      RECT 15.405 1.58 15.765 2.15 ;
      RECT 15.405 0.845 15.575 1.58 ;
      RECT 14.765 0.595 15.575 0.845 ;
      RECT 10.655 2.055 10.985 2.215 ;
      RECT 10.655 1.885 13.015 2.055 ;
      RECT 11.475 2.055 11.805 2.235 ;
    LAYER mcon ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 1.58 15.685 1.75 ;
      RECT 15.515 2.735 15.685 2.905 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 2.735 15.205 2.905 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.24 1.58 10.41 1.75 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 1.58 5.125 1.75 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 19.835 -0.085 20.005 0.085 ;
      RECT 19.835 3.245 20.005 3.415 ;
      RECT 19.355 -0.085 19.525 0.085 ;
      RECT 19.355 3.245 19.525 3.415 ;
      RECT 18.875 -0.085 19.045 0.085 ;
      RECT 18.875 3.245 19.045 3.415 ;
      RECT 18.395 -0.085 18.565 0.085 ;
      RECT 18.395 3.245 18.565 3.415 ;
      RECT 17.915 -0.085 18.085 0.085 ;
      RECT 17.915 3.245 18.085 3.415 ;
      RECT 17.435 -0.085 17.605 0.085 ;
      RECT 17.435 3.245 17.605 3.415 ;
      RECT 16.955 -0.085 17.125 0.085 ;
      RECT 16.955 3.245 17.125 3.415 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 2.735 16.165 2.905 ;
      RECT 15.995 3.245 16.165 3.415 ;
    LAYER met1 ;
      RECT 4.895 1.735 5.185 1.78 ;
      RECT 4.895 1.595 15.745 1.735 ;
      RECT 10.18 1.735 10.47 1.78 ;
      RECT 15.455 1.735 15.745 1.78 ;
      RECT 4.895 1.55 5.185 1.595 ;
      RECT 10.18 1.55 10.47 1.595 ;
      RECT 15.455 1.55 15.745 1.595 ;
  END
END scs8ls_lpflow_srsdfstp_4

MACRO scs8ls_lpflow_srsdfxtp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 13.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.795 1.18 2.275 1.54 ;
        RECT 1.795 1.01 1.965 1.18 ;
        RECT 0.425 0.985 1.965 1.01 ;
        RECT 0.425 1.01 0.755 1.315 ;
        RECT 0.585 0.84 1.965 0.985 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.02 0.255 11.37 0.65 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END SLEEPB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.18 1.59 1.51 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075 1.75 2.49 2.15 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 9.66 1.47 10.56 1.8 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.03 0.345 13.305 1.145 ;
        RECT 13.125 1.145 13.305 1.82 ;
        RECT 12.975 1.82 13.305 2.97 ;
    END
    ANTENNADIFFAREA 0.5673 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.92 3.575 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 13.85 2.945 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 2.735 10.885 2.905 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 2.735 9.925 2.905 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
    LAYER li1 ;
      RECT 12.03 1.645 12.34 2.5 ;
      RECT 12.03 1.315 12.955 1.645 ;
      RECT 12.03 0.42 12.425 1.315 ;
      RECT 8.07 2.435 11.86 2.52 ;
      RECT 6.91 2.35 11.86 2.435 ;
      RECT 11.69 1.795 11.86 2.35 ;
      RECT 11.56 1.47 11.86 1.795 ;
      RECT 8.07 2.52 8.745 2.98 ;
      RECT 6.91 2.435 7.395 2.735 ;
      RECT 6.91 2.265 8.35 2.35 ;
      RECT 6.91 1.595 7.4 2.265 ;
      RECT 6.91 1.425 8.44 1.595 ;
      RECT 8.11 1.595 8.44 1.705 ;
      RECT 6.91 0.925 7.21 1.425 ;
      RECT 6.57 0.595 7.21 0.925 ;
      RECT 0 3.245 13.92 3.415 ;
      RECT 13.475 1.8 13.745 3.245 ;
      RECT 5.41 2.945 5.76 3.245 ;
      RECT 2.4 2.66 2.65 3.245 ;
      RECT 12.53 1.84 12.795 3.245 ;
      RECT 0.565 2.305 0.895 3.245 ;
      RECT 0 -0.085 13.92 0.085 ;
      RECT 13.475 0.085 13.745 1.12 ;
      RECT 11.325 0.935 11.71 1.265 ;
      RECT 11.54 0.085 11.71 0.935 ;
      RECT 12.595 0.085 12.86 1.145 ;
      RECT 2.475 0.085 2.645 0.67 ;
      RECT 4.755 0.085 5.085 0.38 ;
      RECT 7.845 0.085 8.095 0.915 ;
      RECT 0.595 0.085 0.925 0.67 ;
      RECT 10.73 1.99 11.52 2.18 ;
      RECT 10.73 0.99 10.9 1.99 ;
      RECT 10.595 0.82 10.9 0.99 ;
      RECT 10.595 0.765 10.765 0.82 ;
      RECT 8.555 0.585 10.765 0.765 ;
      RECT 8.555 0.765 9.41 0.915 ;
      RECT 10.665 2.69 10.995 3.065 ;
      RECT 8.52 2.095 10.425 2.18 ;
      RECT 7.57 1.985 10.425 2.095 ;
      RECT 9.275 1.285 9.88 1.3 ;
      RECT 9.275 1.13 10.425 1.285 ;
      RECT 9.71 0.955 10.425 1.13 ;
      RECT 7.57 1.875 8.69 1.985 ;
      RECT 9.275 1.3 9.48 1.985 ;
      RECT 7.57 1.765 7.9 1.875 ;
      RECT 9.515 2.69 9.975 3 ;
      RECT 3.16 2.405 3.88 2.735 ;
      RECT 3.16 2.15 3.455 2.405 ;
      RECT 3 1.915 3.455 2.15 ;
      RECT 3 0.69 3.21 1.915 ;
      RECT 2.825 0.505 3.21 0.69 ;
      RECT 2.825 0.425 3.57 0.505 ;
      RECT 2.825 0.255 4.575 0.425 ;
      RECT 4.405 0.425 4.575 0.55 ;
      RECT 4.405 0.55 5.425 0.72 ;
      RECT 5.255 0.425 5.425 0.55 ;
      RECT 5.255 0.255 7.655 0.425 ;
      RECT 6.135 0.425 6.345 1.12 ;
      RECT 7.38 0.425 7.655 1.085 ;
      RECT 6.135 1.12 6.675 1.425 ;
      RECT 7.38 1.085 8.945 1.255 ;
      RECT 8.775 1.255 8.945 1.395 ;
      RECT 8.775 1.395 9.07 1.725 ;
      RECT 4.5 2.77 4.78 2.91 ;
      RECT 4.5 2.6 6.55 2.77 ;
      RECT 6.38 2.77 6.55 2.905 ;
      RECT 4.5 1.895 4.78 2.6 ;
      RECT 6.38 2.905 7.9 3.075 ;
      RECT 3.985 1.725 5.44 1.895 ;
      RECT 7.57 2.745 7.9 2.905 ;
      RECT 5.11 1.23 5.44 1.725 ;
      RECT 3.985 0.675 4.235 1.725 ;
      RECT 5.14 2.105 6.505 2.425 ;
      RECT 5.61 1.06 5.94 2.105 ;
      RECT 4.57 0.89 5.94 1.06 ;
      RECT 4.57 1.06 4.9 1.475 ;
      RECT 5.61 0.595 5.94 0.89 ;
      RECT 1.41 2.32 2.99 2.49 ;
      RECT 2.82 2.49 2.99 2.905 ;
      RECT 2.66 1.18 2.83 2.32 ;
      RECT 2.82 2.905 4.33 3.075 ;
      RECT 2.485 1.01 2.83 1.18 ;
      RECT 4.05 2.235 4.33 2.905 ;
      RECT 2.135 0.84 2.655 1.01 ;
      RECT 3.635 2.065 4.33 2.235 ;
      RECT 2.135 0.67 2.305 0.84 ;
      RECT 3.635 1.005 3.805 2.065 ;
      RECT 1.495 0.5 2.305 0.67 ;
      RECT 3.475 0.675 3.805 1.005 ;
      RECT 1.495 0.34 1.825 0.5 ;
      RECT 1.41 2.49 1.74 3 ;
      RECT 0.085 1.91 1.905 2.08 ;
      RECT 0.585 1.75 1.905 1.91 ;
      RECT 0.085 2.08 0.365 3.045 ;
      RECT 0.085 0.675 0.255 1.91 ;
      RECT 0.085 0.345 0.415 0.675 ;
      RECT 0.585 1.555 0.915 1.75 ;
  END
END scs8ls_lpflow_srsdfxtp_2

MACRO scs8ls_lpflow_srsdfxtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 14.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.795 1.18 2.275 1.54 ;
        RECT 1.795 1.01 1.965 1.18 ;
        RECT 0.425 0.985 1.965 1.01 ;
        RECT 0.425 1.01 0.755 1.315 ;
        RECT 0.585 0.84 1.965 0.985 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.02 0.255 11.37 0.65 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END SLEEPB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.18 1.59 1.51 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075 1.75 2.49 2.15 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 9.66 1.47 10.56 1.8 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.03 0.345 13.305 1.145 ;
        RECT 13.125 1.145 13.305 1.46 ;
        RECT 13.125 1.46 14.175 1.545 ;
        RECT 13.125 1.545 14.25 1.63 ;
        RECT 13.915 0.35 14.175 1.46 ;
        RECT 13.125 1.63 13.305 1.82 ;
        RECT 13.915 1.63 14.25 2.97 ;
        RECT 12.975 1.82 13.305 2.97 ;
    END
    ANTENNADIFFAREA 1.1346 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 14.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 14.88 3.575 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 14.81 2.945 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 2.735 10.885 2.905 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 2.735 9.925 2.905 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
    LAYER li1 ;
      RECT 12.03 1.645 12.34 2.98 ;
      RECT 12.03 1.315 12.955 1.645 ;
      RECT 12.03 0.35 12.425 1.315 ;
      RECT 8.07 2.435 11.86 2.52 ;
      RECT 6.91 2.35 11.86 2.435 ;
      RECT 11.69 1.795 11.86 2.35 ;
      RECT 11.56 1.47 11.86 1.795 ;
      RECT 8.07 2.52 8.745 2.98 ;
      RECT 6.91 2.435 7.395 2.735 ;
      RECT 6.91 2.265 8.35 2.35 ;
      RECT 6.91 1.595 7.4 2.265 ;
      RECT 6.91 1.425 8.44 1.595 ;
      RECT 8.11 1.595 8.44 1.705 ;
      RECT 6.91 0.925 7.21 1.425 ;
      RECT 6.57 0.595 7.21 0.925 ;
      RECT 10.73 1.99 11.52 2.18 ;
      RECT 10.73 0.99 10.9 1.99 ;
      RECT 10.595 0.82 10.9 0.99 ;
      RECT 10.595 0.765 10.765 0.82 ;
      RECT 8.555 0.585 10.765 0.765 ;
      RECT 8.555 0.765 9.41 0.915 ;
      RECT 0 3.245 14.88 3.415 ;
      RECT 14.42 1.8 14.67 3.245 ;
      RECT 5.41 2.945 5.76 3.245 ;
      RECT 2.4 2.66 2.65 3.245 ;
      RECT 12.53 1.84 12.795 3.245 ;
      RECT 13.475 1.8 13.745 3.245 ;
      RECT 0.565 2.305 0.895 3.245 ;
      RECT 0 -0.085 14.88 0.085 ;
      RECT 14.345 0.085 14.63 1.12 ;
      RECT 11.325 0.935 11.71 1.265 ;
      RECT 11.54 0.085 11.71 0.935 ;
      RECT 12.595 0.085 12.86 1.145 ;
      RECT 13.475 0.085 13.745 1.12 ;
      RECT 2.475 0.085 2.645 0.67 ;
      RECT 4.755 0.085 5.085 0.38 ;
      RECT 7.845 0.085 8.095 0.915 ;
      RECT 0.595 0.085 0.925 0.67 ;
      RECT 10.665 2.69 10.995 3.065 ;
      RECT 8.52 2.095 10.425 2.18 ;
      RECT 7.57 1.985 10.425 2.095 ;
      RECT 9.275 1.285 9.88 1.3 ;
      RECT 9.275 1.13 10.425 1.285 ;
      RECT 9.71 0.955 10.425 1.13 ;
      RECT 7.57 1.875 8.69 1.985 ;
      RECT 9.275 1.3 9.48 1.985 ;
      RECT 7.57 1.765 7.9 1.875 ;
      RECT 9.515 2.69 9.975 3 ;
      RECT 3.16 2.405 3.88 2.735 ;
      RECT 3.16 2.15 3.455 2.405 ;
      RECT 3 1.915 3.455 2.15 ;
      RECT 3 0.69 3.21 1.915 ;
      RECT 2.825 0.505 3.21 0.69 ;
      RECT 2.825 0.425 3.57 0.505 ;
      RECT 2.825 0.255 4.575 0.425 ;
      RECT 4.405 0.425 4.575 0.55 ;
      RECT 4.405 0.55 5.425 0.72 ;
      RECT 5.255 0.425 5.425 0.55 ;
      RECT 5.255 0.255 7.655 0.425 ;
      RECT 6.135 0.425 6.345 1.12 ;
      RECT 7.38 0.425 7.655 1.085 ;
      RECT 6.135 1.12 6.675 1.425 ;
      RECT 7.38 1.085 8.945 1.255 ;
      RECT 8.775 1.255 8.945 1.395 ;
      RECT 8.775 1.395 9.07 1.725 ;
      RECT 4.5 2.77 4.78 2.91 ;
      RECT 4.5 2.6 6.55 2.77 ;
      RECT 6.38 2.77 6.55 2.905 ;
      RECT 4.5 1.895 4.78 2.6 ;
      RECT 6.38 2.905 7.9 3.075 ;
      RECT 3.985 1.725 5.44 1.895 ;
      RECT 7.57 2.745 7.9 2.905 ;
      RECT 5.11 1.23 5.44 1.725 ;
      RECT 3.985 0.675 4.235 1.725 ;
      RECT 5.14 2.105 6.505 2.425 ;
      RECT 5.61 1.06 5.94 2.105 ;
      RECT 4.57 0.89 5.94 1.06 ;
      RECT 4.57 1.06 4.9 1.475 ;
      RECT 5.61 0.595 5.94 0.89 ;
      RECT 1.41 2.32 2.99 2.49 ;
      RECT 2.82 2.49 2.99 2.905 ;
      RECT 2.66 1.18 2.83 2.32 ;
      RECT 2.82 2.905 4.33 3.075 ;
      RECT 2.485 1.01 2.83 1.18 ;
      RECT 4.05 2.235 4.33 2.905 ;
      RECT 2.135 0.84 2.655 1.01 ;
      RECT 3.635 2.065 4.33 2.235 ;
      RECT 2.135 0.67 2.305 0.84 ;
      RECT 3.635 1.005 3.805 2.065 ;
      RECT 1.495 0.5 2.305 0.67 ;
      RECT 3.475 0.675 3.805 1.005 ;
      RECT 1.495 0.34 1.825 0.5 ;
      RECT 1.41 2.49 1.74 3 ;
      RECT 0.085 1.91 1.905 2.08 ;
      RECT 0.585 1.75 1.905 1.91 ;
      RECT 0.085 2.08 0.365 3.045 ;
      RECT 0.085 0.675 0.255 1.91 ;
      RECT 0.085 0.345 0.415 0.675 ;
      RECT 0.585 1.555 0.915 1.75 ;
  END
END scs8ls_lpflow_srsdfxtp_4

MACRO scs8ls_lpflow_sleep_pargate
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 8.64 BY 3.33 ;
  SYMMETRY X Y R90 ;
  SITE unit ;

  PIN sleep
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.105 0.41 8.53 2.92 ;
    END
    ANTENNAGATEAREA 7.56 ;
  END sleep

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 8.64 0.245 ;
    END
  END vgnd

  PIN realvpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 0.805 0 1.595 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 6.285 0 7.055 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.465 0 5.235 3.33 ;
    END
    PORT
      LAYER met2 ;
        RECT 2.645 0 3.415 3.33 ;
    END
    PORT
      LAYER via ;
        RECT 4.52 2.33 4.67 2.48 ;
        RECT 4.55 0.78 4.7 0.93 ;
        RECT 5.03 2.33 5.18 2.48 ;
        RECT 5 0.78 5.15 0.93 ;
        RECT 6.37 0.78 6.52 0.93 ;
        RECT 6.34 2.33 6.49 2.48 ;
        RECT 6.82 0.78 6.97 0.93 ;
        RECT 6.82 2.33 6.97 2.48 ;
        RECT 3.18 0.78 3.33 0.93 ;
        RECT 3.21 2.33 3.36 2.48 ;
        RECT 2.73 0.78 2.88 0.93 ;
        RECT 2.7 2.33 2.85 2.48 ;
        RECT 1.36 0.78 1.51 0.93 ;
        RECT 1.39 2.33 1.54 2.48 ;
        RECT 0.89 0.78 1.04 0.93 ;
        RECT 0.89 2.33 1.04 2.48 ;
    END
  END realvpwr

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 1.735 0 2.505 3.49 ;
    END
    PORT
      LAYER met2 ;
        RECT 7.195 0 7.965 3.49 ;
    END
    PORT
      LAYER met2 ;
        RECT 5.375 0 6.145 3.49 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.555 0 4.325 3.49 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 3.085 8.64 3.575 ;
    END
    PORT
      LAYER via ;
        RECT 4.09 0.44 4.24 0.59 ;
        RECT 7.25 3.255 7.4 3.405 ;
        RECT 3.64 0.44 3.79 0.59 ;
        RECT 4.12 3.255 4.27 3.405 ;
        RECT 7.76 3.255 7.91 3.405 ;
        RECT 7.73 0.44 7.88 0.59 ;
        RECT 5.91 0.44 6.06 0.59 ;
        RECT 5.43 3.255 5.58 3.405 ;
        RECT 5.46 0.44 5.61 0.59 ;
        RECT 5.94 3.255 6.09 3.405 ;
        RECT 2.27 0.44 2.42 0.59 ;
        RECT 3.61 3.255 3.76 3.405 ;
        RECT 2.3 3.255 2.45 3.405 ;
        RECT 1.82 0.44 1.97 0.59 ;
        RECT 1.79 3.255 1.94 3.405 ;
        RECT 7.28 0.44 7.43 0.59 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 0.805 2.275 7.055 2.535 ;
      RECT 0.805 0.785 7.055 0.985 ;
      RECT 0.805 0.725 1.595 0.785 ;
      RECT 2.645 0.725 3.415 0.785 ;
      RECT 4.465 0.725 5.235 0.785 ;
      RECT 6.285 0.725 7.055 0.785 ;
      RECT 1.735 0.585 2.505 0.645 ;
      RECT 1.735 0.385 7.965 0.585 ;
      RECT 3.555 0.585 4.325 0.645 ;
      RECT 5.375 0.585 6.145 0.645 ;
      RECT 7.195 0.585 7.965 0.645 ;
    LAYER li1 ;
      RECT 0 3.245 8.64 3.415 ;
      RECT 0.775 2.9 7.935 3.245 ;
      RECT 1.75 1.95 2.495 2.9 ;
      RECT 3.57 1.95 4.305 2.9 ;
      RECT 5.385 1.95 6.13 2.9 ;
      RECT 7.185 1.95 7.935 2.9 ;
      RECT 0.945 1.78 1.58 2.73 ;
      RECT 0.775 1.55 7.855 1.78 ;
      RECT 2.665 1.78 3.4 2.73 ;
      RECT 4.475 1.78 5.215 2.73 ;
      RECT 6.3 1.78 7.015 2.73 ;
      RECT 0.945 0.6 1.58 1.55 ;
      RECT 2.665 0.6 3.4 1.55 ;
      RECT 4.475 0.6 5.215 1.55 ;
      RECT 6.3 0.6 7.015 1.55 ;
      RECT 1.75 0.43 2.495 1.38 ;
      RECT 0.775 0.2 7.935 0.43 ;
      RECT 3.57 0.43 4.305 1.38 ;
      RECT 5.385 0.43 6.13 1.38 ;
      RECT 7.185 0.43 7.935 1.38 ;
    LAYER mcon ;
      RECT 6.815 0.77 6.985 0.94 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 7.255 0.43 7.425 0.6 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.735 0.43 7.905 0.6 ;
      RECT 5.435 0.43 5.605 0.6 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 5.005 0.77 5.175 0.94 ;
      RECT 5.015 2.32 5.185 2.49 ;
      RECT 4.525 0.77 4.695 0.94 ;
      RECT 4.505 2.32 4.675 2.49 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 4.095 0.43 4.265 0.6 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 3.615 0.43 3.785 0.6 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 3.185 0.77 3.355 0.94 ;
      RECT 3.2 2.32 3.37 2.49 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 2.705 0.77 2.875 0.94 ;
      RECT 2.695 2.32 2.865 2.49 ;
      RECT 2.275 0.43 2.445 0.6 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.795 0.43 1.965 0.6 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.365 0.77 1.535 0.94 ;
      RECT 1.38 2.32 1.55 2.49 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.945 0.77 1.115 0.94 ;
      RECT 0.945 2.32 1.115 2.49 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 6.33 2.32 6.5 2.49 ;
      RECT 6.345 0.77 6.515 0.94 ;
      RECT 6.815 2.32 6.985 2.49 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 5.915 0.43 6.085 0.6 ;
  END
END scs8ls_lpflow_sleep_pargate

MACRO scs8ls_lpflow_srsdfrtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 20.64 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 20.205 0.35 20.535 1.82 ;
        RECT 19.995 1.82 20.535 2.155 ;
        RECT 19.995 2.155 20.325 2.975 ;
    END
    ANTENNADIFFAREA 0.5395 ;
  END Q

  PIN RESETB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.92 1.55 4.25 1.88 ;
    END
    ANTENNAGATEAREA 0.598 ;
  END RESETB

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.5 0.935 2.17 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.84 2.135 2.17 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.35 1.55 3.715 1.88 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 16.59 1.46 17.155 1.79 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END CLK

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.235 1.12 18.565 1.45 ;
    END
    ANTENNAGATEAREA 0.598 ;
  END SLEEPB

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 20.64 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 20.64 3.575 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 20.57 2.945 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 15.035 2.735 15.205 2.905 ;
      RECT 15.515 2.735 15.685 2.905 ;
      RECT 17.435 2.735 17.605 2.905 ;
      RECT 15.995 2.735 16.165 2.905 ;
      RECT 20.315 -0.085 20.485 0.085 ;
      RECT 20.315 3.245 20.485 3.415 ;
      RECT 19.835 -0.085 20.005 0.085 ;
      RECT 19.835 3.245 20.005 3.415 ;
      RECT 19.355 -0.085 19.525 0.085 ;
      RECT 19.355 3.245 19.525 3.415 ;
      RECT 18.875 -0.085 19.045 0.085 ;
      RECT 18.875 3.245 19.045 3.415 ;
      RECT 18.395 -0.085 18.565 0.085 ;
      RECT 18.395 3.245 18.565 3.415 ;
      RECT 17.915 -0.085 18.085 0.085 ;
      RECT 17.915 3.245 18.085 3.415 ;
      RECT 17.435 -0.085 17.605 0.085 ;
      RECT 17.435 3.245 17.605 3.415 ;
      RECT 16.955 -0.085 17.125 0.085 ;
      RECT 16.955 2.735 17.125 2.905 ;
      RECT 16.955 3.245 17.125 3.415 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 16.475 2.735 16.645 2.905 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 2.735 14.725 2.905 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
    LAYER li1 ;
      RECT 12.21 2.35 19.325 2.52 ;
      RECT 19.155 1.645 19.325 2.35 ;
      RECT 19.075 1.315 19.345 1.645 ;
      RECT 9.835 2.565 12.54 2.735 ;
      RECT 12.21 2.52 12.54 2.565 ;
      RECT 9.835 2.04 10.5 2.565 ;
      RECT 10.19 0.605 10.5 2.04 ;
      RECT 13.625 2.52 13.955 2.97 ;
      RECT 16.25 1.74 16.42 2.35 ;
      RECT 15.985 1.41 16.42 1.74 ;
      RECT 17.895 1.85 18.49 2.18 ;
      RECT 16.93 0.78 18.345 0.95 ;
      RECT 18.015 0.345 18.345 0.78 ;
      RECT 17.895 0.95 18.065 1.85 ;
      RECT 16.93 0.425 17.1 0.78 ;
      RECT 14.985 0.255 17.1 0.425 ;
      RECT 14.985 0.425 15.315 0.6 ;
      RECT 14.015 0.6 15.315 0.77 ;
      RECT 14.015 0.77 14.185 1.32 ;
      RECT 12.93 1.32 14.185 1.5 ;
      RECT 16.855 2.01 17.495 2.18 ;
      RECT 17.325 1.29 17.495 2.01 ;
      RECT 16.59 1.12 17.495 1.29 ;
      RECT 16.105 1.11 16.76 1.12 ;
      RECT 14.355 0.95 16.76 1.11 ;
      RECT 14.355 1.11 14.525 1.67 ;
      RECT 14.355 0.94 16.435 0.95 ;
      RECT 11.64 1.67 14.525 1.84 ;
      RECT 16.105 0.595 16.435 0.94 ;
      RECT 11.64 1.51 11.97 1.67 ;
      RECT 11.1 2.01 16.08 2.18 ;
      RECT 14.695 1.93 16.08 2.01 ;
      RECT 11.1 1.325 11.43 2.01 ;
      RECT 14.695 1.28 14.955 1.93 ;
      RECT 11.1 1.155 12.235 1.325 ;
      RECT 11.905 0.575 12.235 1.155 ;
      RECT 14.525 2.69 17.73 3.025 ;
      RECT 12.695 0.98 13.845 1.15 ;
      RECT 12.695 0.575 12.945 0.98 ;
      RECT 13.675 0.575 13.845 0.98 ;
      RECT 8.555 2.905 13.455 3.075 ;
      RECT 8.555 2.825 8.725 2.905 ;
      RECT 13.125 2.745 13.455 2.905 ;
      RECT 8.395 2.435 8.725 2.825 ;
      RECT 5.78 2.43 8.725 2.435 ;
      RECT 5.78 2.435 7.68 2.6 ;
      RECT 7.51 2.265 8.725 2.43 ;
      RECT 4.925 2.6 5.95 2.77 ;
      RECT 8.395 1.665 8.725 2.265 ;
      RECT 4.925 1.92 5.095 2.6 ;
      RECT 8.395 1.495 9.4 1.665 ;
      RECT 4.885 1.59 5.215 1.92 ;
      RECT 9.07 1.665 9.4 1.825 ;
      RECT 8.395 1.335 8.99 1.495 ;
      RECT 7.32 1.845 8.135 2.095 ;
      RECT 7.965 1.175 8.135 1.845 ;
      RECT 6.28 1.165 8.135 1.175 ;
      RECT 6.28 1.175 6.61 1.485 ;
      RECT 6.28 1.005 9.53 1.165 ;
      RECT 9.2 1.165 9.53 1.285 ;
      RECT 7.59 0.995 9.53 1.005 ;
      RECT 7.59 0.575 7.84 0.995 ;
      RECT 9.2 0.435 9.53 0.995 ;
      RECT 9.2 0.265 10.93 0.435 ;
      RECT 10.68 0.435 10.93 2.395 ;
      RECT 5.265 2.26 5.555 2.43 ;
      RECT 5.265 2.09 7.11 2.26 ;
      RECT 6.78 1.675 7.11 2.09 ;
      RECT 5.385 1.265 5.555 2.09 ;
      RECT 6.78 1.345 7.795 1.675 ;
      RECT 5.375 0.935 5.555 1.265 ;
      RECT 4.615 0.425 4.865 1.08 ;
      RECT 4.615 0.255 6.59 0.425 ;
      RECT 6.26 0.425 6.59 0.835 ;
      RECT 2.305 2.1 4.755 2.24 ;
      RECT 4.47 2.24 4.755 2.99 ;
      RECT 2.98 2.07 4.715 2.1 ;
      RECT 4.545 1.42 4.715 2.07 ;
      RECT 4.545 1.25 5.205 1.42 ;
      RECT 5.035 0.765 5.205 1.25 ;
      RECT 5.035 0.595 6.055 0.765 ;
      RECT 5.725 0.765 6.055 1.265 ;
      RECT 1.96 2.51 2.635 2.99 ;
      RECT 1.225 2.34 2.635 2.51 ;
      RECT 2.305 2.325 2.635 2.34 ;
      RECT 2.305 2.24 3.08 2.325 ;
      RECT 1.225 1.5 2.08 1.67 ;
      RECT 1.83 0.935 2.08 1.5 ;
      RECT 1.225 1.67 1.395 2.34 ;
      RECT 2.645 1.21 4.375 1.38 ;
      RECT 2.645 0.74 2.975 1.21 ;
      RECT 4.045 0.58 4.375 1.21 ;
      RECT 1.07 0.425 1.32 0.99 ;
      RECT 1.07 0.255 3.405 0.425 ;
      RECT 3.155 0.425 3.405 1.04 ;
      RECT 2.305 1.6 2.88 1.93 ;
      RECT 2.305 0.765 2.475 1.6 ;
      RECT 1.49 0.595 2.475 0.765 ;
      RECT 1.49 0.765 1.66 1.16 ;
      RECT 0.105 1.16 1.66 1.33 ;
      RECT 0.105 1.33 0.435 2.99 ;
      RECT 0.105 0.53 0.355 1.16 ;
      RECT 0 -0.085 20.64 0.085 ;
      RECT 18.805 0.085 19.055 0.805 ;
      RECT 19.855 0.085 20.025 1.13 ;
      RECT 0.535 0.085 0.865 0.99 ;
      RECT 3.615 0.085 3.865 1.04 ;
      RECT 7.05 0.085 7.38 0.835 ;
      RECT 8.02 0.085 8.35 0.825 ;
      RECT 11.365 0.085 11.695 0.985 ;
      RECT 13.125 0.085 13.455 0.81 ;
      RECT 17.475 0.085 17.805 0.61 ;
      RECT 0 3.245 20.64 3.415 ;
      RECT 6.12 2.77 6.45 3.245 ;
      RECT 7.85 2.605 8.18 3.245 ;
      RECT 3.245 2.41 4.3 3.245 ;
      RECT 19.495 1.815 19.825 3.245 ;
      RECT 0.645 2.34 0.975 3.245 ;
      RECT 19.515 1.315 20.02 1.645 ;
      RECT 18.735 1.815 18.985 2.18 ;
      RECT 18.735 1.145 18.905 1.815 ;
      RECT 18.735 0.975 19.685 1.145 ;
      RECT 19.515 1.145 19.685 1.315 ;
      RECT 19.235 0.345 19.685 0.975 ;
  END
END scs8ls_lpflow_srsdfrtp_1

MACRO scs8ls_lpflow_srsdfstp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 18.72 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SETB
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.725 0.78 7.16 1.03 ;
        RECT 6.725 1.03 7.22 1.265 ;
    END
    ANTENNAGATEAREA 0.439 ;
  END SETB

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.365 0.35 18.62 3.075 ;
    END
    ANTENNADIFFAREA 0.519 ;
  END Q

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.545 1.43 1.875 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.725 1.18 3.235 1.555 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.205 0.835 1.875 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.935 1.22 16.26 2.15 ;
    END
    ANTENNAGATEAREA 0.598 ;
  END SLEEPB

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 14.965 1.18 15.235 2.15 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END CLK

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 18.72 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 18.72 3.575 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 18.65 2.945 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 15.515 2.735 15.685 2.905 ;
      RECT 18.395 -0.085 18.565 0.085 ;
      RECT 18.395 3.245 18.565 3.415 ;
      RECT 17.915 -0.085 18.085 0.085 ;
      RECT 17.915 3.245 18.085 3.415 ;
      RECT 17.435 -0.085 17.605 0.085 ;
      RECT 17.435 3.245 17.605 3.415 ;
      RECT 16.955 -0.085 17.125 0.085 ;
      RECT 16.955 3.245 17.125 3.415 ;
      RECT 16.475 -0.085 16.645 0.085 ;
      RECT 16.475 3.245 16.645 3.415 ;
      RECT 15.995 -0.085 16.165 0.085 ;
      RECT 15.995 2.735 16.165 2.905 ;
      RECT 15.995 3.245 16.165 3.415 ;
      RECT 15.515 -0.085 15.685 0.085 ;
      RECT 15.515 1.58 15.685 1.75 ;
      RECT 15.515 3.245 15.685 3.415 ;
      RECT 15.035 -0.085 15.205 0.085 ;
      RECT 15.035 2.735 15.205 2.905 ;
      RECT 15.035 3.245 15.205 3.415 ;
      RECT 14.555 -0.085 14.725 0.085 ;
      RECT 14.555 3.245 14.725 3.415 ;
      RECT 14.075 -0.085 14.245 0.085 ;
      RECT 14.075 3.245 14.245 3.415 ;
      RECT 13.595 -0.085 13.765 0.085 ;
      RECT 13.595 3.245 13.765 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.24 1.58 10.41 1.75 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 1.58 5.125 1.75 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
    LAYER met1 ;
      RECT 4.895 1.735 5.185 1.78 ;
      RECT 4.895 1.595 15.745 1.735 ;
      RECT 10.18 1.735 10.47 1.78 ;
      RECT 15.455 1.735 15.745 1.78 ;
      RECT 4.895 1.55 5.185 1.595 ;
      RECT 10.18 1.55 10.47 1.595 ;
      RECT 15.455 1.55 15.745 1.595 ;
    LAYER li1 ;
      RECT 15.405 1.58 15.765 2.15 ;
      RECT 15.405 0.845 15.575 1.58 ;
      RECT 14.765 0.595 15.575 0.845 ;
      RECT 10.655 2.055 10.985 2.215 ;
      RECT 10.655 1.885 13.015 2.055 ;
      RECT 11.475 2.055 11.805 2.235 ;
      RECT 12.845 1.055 13.015 1.885 ;
      RECT 12.845 0.885 14.55 1.055 ;
      RECT 14.22 1.055 14.55 1.26 ;
      RECT 7.845 2.905 8.695 3.075 ;
      RECT 8.525 1.74 8.695 2.905 ;
      RECT 7.845 1.605 8.015 2.905 ;
      RECT 8.525 1.355 8.755 1.74 ;
      RECT 5.65 1.45 8.015 1.605 ;
      RECT 8.525 0.765 8.695 1.355 ;
      RECT 5.65 1.605 6.895 1.62 ;
      RECT 6.725 1.435 8.015 1.45 ;
      RECT 8.525 0.595 9.535 0.765 ;
      RECT 7.845 1.37 8.015 1.435 ;
      RECT 9.365 0.765 9.535 2.405 ;
      RECT 9.365 2.405 12.145 2.575 ;
      RECT 11.975 2.395 12.145 2.405 ;
      RECT 11.975 2.225 13.355 2.395 ;
      RECT 13.185 2.18 13.355 2.225 ;
      RECT 13.185 2.01 14.21 2.18 ;
      RECT 14.04 1.8 14.21 2.01 ;
      RECT 14.04 1.55 14.37 1.8 ;
      RECT 5.65 0.92 5.82 1.45 ;
      RECT 5.08 0.75 5.82 0.92 ;
      RECT 5.08 0.425 5.25 0.75 ;
      RECT 3.42 0.255 5.25 0.425 ;
      RECT 3.42 0.425 4.015 0.555 ;
      RECT 3.42 0.555 3.67 1.695 ;
      RECT 3.42 1.695 4.255 2.025 ;
      RECT 4.005 2.025 4.255 2.395 ;
      RECT 10.425 1.205 11.455 1.375 ;
      RECT 10.425 0.605 10.595 1.205 ;
      RECT 11.205 0.605 11.455 1.205 ;
      RECT 10.165 1.545 10.415 2.145 ;
      RECT 8.185 1.2 8.355 2.565 ;
      RECT 7.825 0.595 8.355 1.2 ;
      RECT 6.68 2.485 7.01 2.58 ;
      RECT 5.9 2.29 7.01 2.485 ;
      RECT 5.9 2.13 6.23 2.29 ;
      RECT 5.31 1.79 6.77 1.96 ;
      RECT 6.44 1.96 6.77 2.015 ;
      RECT 5.205 2.67 5.535 3 ;
      RECT 5.31 1.96 5.48 2.67 ;
      RECT 5.31 1.26 5.48 1.79 ;
      RECT 4.745 1.135 5.48 1.26 ;
      RECT 4.41 1.09 5.48 1.135 ;
      RECT 4.41 0.82 4.91 1.09 ;
      RECT 5.99 1.09 6.555 1.27 ;
      RECT 6.305 0.595 6.555 1.09 ;
      RECT 4.77 1.58 5.125 2.035 ;
      RECT 3.665 2.655 5.035 2.825 ;
      RECT 3.665 2.395 3.835 2.655 ;
      RECT 4.43 1.525 4.6 2.655 ;
      RECT 1.44 2.225 3.835 2.395 ;
      RECT 3.98 1.355 4.6 1.525 ;
      RECT 3.98 0.755 4.23 1.355 ;
      RECT 1.44 2.395 1.77 2.735 ;
      RECT 1.6 1.035 1.77 2.225 ;
      RECT 0.92 0.865 1.77 1.035 ;
      RECT 0.92 0.575 1.25 0.865 ;
      RECT 1.94 1.725 2.74 2.055 ;
      RECT 2.385 0.675 2.74 1.01 ;
      RECT 1.94 1.305 2.555 1.725 ;
      RECT 2.385 1.01 2.555 1.305 ;
      RECT 1.02 2.905 2.22 3.075 ;
      RECT 1.97 2.65 2.22 2.905 ;
      RECT 1.02 2.215 1.19 2.905 ;
      RECT 0.1 2.045 1.19 2.215 ;
      RECT 0.1 2.215 0.43 3.065 ;
      RECT 0 -0.085 18.72 0.085 ;
      RECT 7.33 0.085 7.5 0.895 ;
      RECT 10.775 0.085 11.025 1.035 ;
      RECT 11.745 0.085 11.995 0.955 ;
      RECT 16.085 0.085 16.335 0.71 ;
      RECT 17.86 0.085 18.19 1.015 ;
      RECT 0.1 0.085 0.43 1.035 ;
      RECT 1.94 0.085 2.19 1.035 ;
      RECT 2.92 0.085 3.25 1.01 ;
      RECT 5.465 0.085 5.795 0.58 ;
      RECT 0 3.245 18.72 3.415 ;
      RECT 17.855 1.815 18.185 3.245 ;
      RECT 6.085 2.75 6.415 3.245 ;
      RECT 2.925 2.565 3.255 3.245 ;
      RECT 7.25 2.29 7.58 3.245 ;
      RECT 0.6 2.385 0.85 3.245 ;
      RECT 17.39 1.995 17.675 2.675 ;
      RECT 17.505 1.55 17.675 1.995 ;
      RECT 17.505 1.22 18.18 1.55 ;
      RECT 17.505 0.675 17.675 1.22 ;
      RECT 17.325 0.35 17.675 0.675 ;
      RECT 13.8 2.35 17.22 2.49 ;
      RECT 14.425 2.32 17.22 2.35 ;
      RECT 17.05 1.825 17.22 2.32 ;
      RECT 17.005 1.495 17.335 1.825 ;
      RECT 8.925 2.745 12.485 3.075 ;
      RECT 12.315 2.735 12.485 2.745 ;
      RECT 8.925 2.235 9.195 2.745 ;
      RECT 12.315 2.565 14.13 2.735 ;
      RECT 8.925 1.225 9.095 2.235 ;
      RECT 13.8 2.52 14.13 2.565 ;
      RECT 8.865 0.935 9.195 1.225 ;
      RECT 13.8 2.49 14.595 2.52 ;
      RECT 15.745 0.88 16.835 1.05 ;
      RECT 16.455 1.05 16.835 2.15 ;
      RECT 16.665 0.8 16.835 0.88 ;
      RECT 16.665 0.63 17.125 0.8 ;
      RECT 16.795 0.42 17.125 0.63 ;
      RECT 12.165 0.255 15.915 0.425 ;
      RECT 15.745 0.425 15.915 0.88 ;
      RECT 11.625 1.125 12.335 1.375 ;
      RECT 12.165 0.425 12.335 1.125 ;
      RECT 13.32 0.425 13.65 0.715 ;
      RECT 12.655 2.905 16.305 3.075 ;
      RECT 14.905 2.66 16.305 2.905 ;
  END
END scs8ls_lpflow_srsdfstp_1

MACRO scs8ls_lpflow_srsdfxtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 13.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.795 1.18 2.275 1.54 ;
        RECT 1.795 1.01 1.965 1.18 ;
        RECT 0.425 0.985 1.965 1.01 ;
        RECT 0.425 1.01 0.755 1.315 ;
        RECT 0.585 0.84 1.965 0.985 ;
    END
    ANTENNAGATEAREA 0.318 ;
  END SCE

  PIN SLEEPB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.02 0.255 11.37 0.65 ;
    END
    ANTENNAGATEAREA 0.222 ;
  END SLEEPB

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.18 1.59 1.51 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END D

  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075 1.75 2.49 2.15 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END SCD

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 9.66 1.47 10.56 1.8 ;
    END
    ANTENNAGATEAREA 0.159 ;
  END CLK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.03 0.345 13.305 1.145 ;
        RECT 13.125 1.145 13.305 1.82 ;
        RECT 12.975 1.82 13.305 2.97 ;
    END
    ANTENNADIFFAREA 0.5041 ;
  END Q

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 13.44 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 13.44 3.575 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 13.37 2.945 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 13.115 -0.085 13.285 0.085 ;
      RECT 13.115 3.245 13.285 3.415 ;
      RECT 12.635 -0.085 12.805 0.085 ;
      RECT 12.635 3.245 12.805 3.415 ;
      RECT 12.155 -0.085 12.325 0.085 ;
      RECT 12.155 3.245 12.325 3.415 ;
      RECT 11.675 -0.085 11.845 0.085 ;
      RECT 11.675 3.245 11.845 3.415 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 2.735 10.885 2.905 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 2.735 9.925 2.905 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
    LAYER li1 ;
      RECT 10.665 2.69 10.995 3.065 ;
      RECT 8.52 2.095 10.425 2.18 ;
      RECT 7.57 1.985 10.425 2.095 ;
      RECT 9.275 1.285 9.88 1.3 ;
      RECT 9.275 1.13 10.425 1.285 ;
      RECT 9.71 0.955 10.425 1.13 ;
      RECT 7.57 1.875 8.69 1.985 ;
      RECT 9.275 1.3 9.48 1.985 ;
      RECT 7.57 1.765 7.9 1.875 ;
      RECT 9.515 2.69 9.975 3 ;
      RECT 3.16 2.405 3.88 2.735 ;
      RECT 3.16 2.15 3.455 2.405 ;
      RECT 3 1.915 3.455 2.15 ;
      RECT 3 0.69 3.21 1.915 ;
      RECT 2.825 0.505 3.21 0.69 ;
      RECT 2.825 0.425 3.57 0.505 ;
      RECT 2.825 0.255 4.575 0.425 ;
      RECT 4.405 0.425 4.575 0.55 ;
      RECT 4.405 0.55 5.425 0.72 ;
      RECT 5.255 0.425 5.425 0.55 ;
      RECT 5.255 0.255 7.655 0.425 ;
      RECT 6.135 0.425 6.345 1.12 ;
      RECT 7.38 0.425 7.655 1.085 ;
      RECT 6.135 1.12 6.675 1.425 ;
      RECT 7.38 1.085 8.945 1.255 ;
      RECT 8.775 1.255 8.945 1.395 ;
      RECT 8.775 1.395 9.07 1.725 ;
      RECT 4.5 2.77 4.78 2.91 ;
      RECT 4.5 2.6 6.55 2.77 ;
      RECT 6.38 2.77 6.55 2.905 ;
      RECT 4.5 1.895 4.78 2.6 ;
      RECT 6.38 2.905 7.9 3.075 ;
      RECT 3.985 1.725 5.44 1.895 ;
      RECT 7.57 2.745 7.9 2.905 ;
      RECT 5.11 1.23 5.44 1.725 ;
      RECT 3.985 0.675 4.235 1.725 ;
      RECT 5.14 2.105 6.505 2.425 ;
      RECT 5.61 1.06 5.94 2.105 ;
      RECT 4.57 0.89 5.94 1.06 ;
      RECT 4.57 1.06 4.9 1.475 ;
      RECT 5.61 0.595 5.94 0.89 ;
      RECT 1.41 2.32 2.99 2.49 ;
      RECT 2.82 2.49 2.99 2.905 ;
      RECT 2.66 1.18 2.83 2.32 ;
      RECT 2.82 2.905 4.33 3.075 ;
      RECT 2.485 1.01 2.83 1.18 ;
      RECT 4.05 2.235 4.33 2.905 ;
      RECT 2.135 0.84 2.655 1.01 ;
      RECT 3.635 2.065 4.33 2.235 ;
      RECT 2.135 0.67 2.305 0.84 ;
      RECT 3.635 1.005 3.805 2.065 ;
      RECT 1.495 0.5 2.305 0.67 ;
      RECT 3.475 0.675 3.805 1.005 ;
      RECT 1.495 0.34 1.825 0.5 ;
      RECT 1.41 2.49 1.74 3 ;
      RECT 0.085 1.91 1.905 2.08 ;
      RECT 0.585 1.75 1.905 1.91 ;
      RECT 0.085 2.08 0.365 3.045 ;
      RECT 0.085 0.675 0.255 1.91 ;
      RECT 0.085 0.345 0.415 0.675 ;
      RECT 0.585 1.555 0.915 1.75 ;
      RECT 8.07 2.435 11.86 2.52 ;
      RECT 6.91 2.35 11.86 2.435 ;
      RECT 11.69 1.795 11.86 2.35 ;
      RECT 11.56 1.47 11.86 1.795 ;
      RECT 8.07 2.52 8.745 2.98 ;
      RECT 6.91 2.435 7.395 2.735 ;
      RECT 6.91 2.265 8.35 2.35 ;
      RECT 6.91 1.595 7.4 2.265 ;
      RECT 6.91 1.425 8.44 1.595 ;
      RECT 8.11 1.595 8.44 1.705 ;
      RECT 6.91 0.925 7.21 1.425 ;
      RECT 6.57 0.595 7.21 0.925 ;
      RECT 12.03 1.645 12.34 2.5 ;
      RECT 12.03 1.315 12.955 1.645 ;
      RECT 12.03 0.42 12.425 1.315 ;
      RECT 0 3.245 13.44 3.415 ;
      RECT 5.41 2.945 5.76 3.245 ;
      RECT 2.4 2.66 2.65 3.245 ;
      RECT 12.53 1.84 12.795 3.245 ;
      RECT 0.565 2.305 0.895 3.245 ;
      RECT 0 -0.085 13.44 0.085 ;
      RECT 11.325 0.935 11.71 1.265 ;
      RECT 11.54 0.085 11.71 0.935 ;
      RECT 12.595 0.085 12.86 1.145 ;
      RECT 2.475 0.085 2.645 0.67 ;
      RECT 4.755 0.085 5.085 0.38 ;
      RECT 7.845 0.085 8.095 0.915 ;
      RECT 0.595 0.085 0.925 0.67 ;
      RECT 10.73 1.99 11.52 2.18 ;
      RECT 10.73 0.99 10.9 1.99 ;
      RECT 10.595 0.82 10.9 0.99 ;
      RECT 10.595 0.765 10.765 0.82 ;
      RECT 8.555 0.585 10.765 0.765 ;
      RECT 8.555 0.765 9.41 0.915 ;
  END
END scs8ls_lpflow_srsdfxtp_1

MACRO scs8ls_lpflow_clkbufkapwr_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475 0.35 1.805 0.79 ;
        RECT 1.565 0.79 1.805 1.82 ;
        RECT 1.345 1.82 1.805 2.98 ;
    END
    ANTENNADIFFAREA 0.4494 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.3 0.835 1.78 ;
    END
    ANTENNAGATEAREA 0.231 ;
  END A

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 1.85 2.945 ;
    END
  END kapwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.845 2.29 1.175 2.98 ;
      RECT 1.005 1.13 1.395 1.63 ;
      RECT 0.115 0.96 1.395 1.13 ;
      RECT 0.345 2.12 0.675 2.98 ;
      RECT 0.345 1.95 1.175 2.12 ;
      RECT 1.005 1.63 1.175 1.95 ;
      RECT 0.115 0.35 0.445 0.96 ;
      RECT 0 -0.085 1.92 0.085 ;
      RECT 0.615 0.085 1.305 0.68 ;
      RECT 0 3.245 1.92 3.415 ;
    LAYER mcon ;
      RECT 0.93 2.715 1.1 2.885 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_clkbufkapwr_1

MACRO scs8ls_lpflow_clkbufkapwr_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.795 1.78 ;
    END
    ANTENNAGATEAREA 0.924 ;
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2.43 1.92 9.01 2.15 ;
    END
    ANTENNADIFFAREA 3.6288 ;
  END X

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 9.53 2.945 ;
    END
  END kapwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 9.6 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 9.6 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER met1 ;
      RECT 2.015 1.18 8.54 1.41 ;
    LAYER li1 ;
      RECT 8.25 1.19 8.545 1.52 ;
      RECT 7.31 1.19 7.63 1.52 ;
      RECT 6.43 1.19 6.73 1.52 ;
      RECT 5.525 1.19 5.83 1.52 ;
      RECT 4.635 1.19 4.94 1.52 ;
      RECT 3.715 1.19 4.035 1.52 ;
      RECT 2.865 1.19 3.145 1.52 ;
      RECT 9.17 1.82 9.48 2.98 ;
      RECT 0 3.245 9.6 3.415 ;
      RECT 0.115 0.085 0.365 0.81 ;
      RECT 0 -0.085 9.6 0.085 ;
      RECT 0.975 0.085 1.225 0.81 ;
      RECT 1.855 0.085 2.185 0.81 ;
      RECT 2.855 0.085 3.065 0.745 ;
      RECT 3.7 0.085 3.935 0.745 ;
      RECT 4.615 0.085 4.88 0.745 ;
      RECT 5.53 0.085 5.805 0.745 ;
      RECT 6.435 0.085 6.715 0.745 ;
      RECT 7.31 0.085 7.645 0.745 ;
      RECT 8.25 0.085 8.555 0.745 ;
      RECT 9.165 0.085 9.485 0.745 ;
      RECT 0.57 2.12 0.9 2.98 ;
      RECT 0.57 1.95 2.135 2.12 ;
      RECT 1.47 2.12 1.8 2.98 ;
      RECT 1.965 1.46 2.135 1.95 ;
      RECT 1.965 1.15 2.29 1.46 ;
      RECT 0.545 1.13 2.29 1.15 ;
      RECT 0.545 0.98 2.135 1.13 ;
      RECT 0.545 0.395 0.795 0.98 ;
      RECT 1.425 0.395 1.675 0.98 ;
      RECT 2 2.29 2.25 2.98 ;
      RECT 6.445 1.82 6.715 2.98 ;
      RECT 6.905 0.395 7.13 2.98 ;
      RECT 7.33 1.82 7.65 2.98 ;
      RECT 7.83 0.395 8.07 2.98 ;
      RECT 8.25 1.82 8.545 2.98 ;
      RECT 8.725 0.395 8.975 2.98 ;
      RECT 2.865 1.82 3.135 2.98 ;
      RECT 3.325 0.745 3.53 2.98 ;
      RECT 3.245 0.395 3.53 0.745 ;
      RECT 3.73 1.82 4.03 2.98 ;
      RECT 4.215 0.745 4.445 2.98 ;
      RECT 4.115 0.395 4.445 0.745 ;
      RECT 4.63 1.82 4.925 2.98 ;
      RECT 5.12 0.745 5.345 2.98 ;
      RECT 5.05 0.395 5.345 0.745 ;
      RECT 5.545 1.82 5.84 2.98 ;
      RECT 6.02 0.745 6.25 2.98 ;
      RECT 5.975 0.395 6.25 0.745 ;
      RECT 1.1 2.29 1.27 2.98 ;
      RECT 2.46 0.745 2.685 2.98 ;
      RECT 2.4 0.395 2.685 0.745 ;
      RECT 0.12 1.95 0.37 2.98 ;
    LAYER mcon ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.1 2.715 1.27 2.885 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 2.715 0.325 2.885 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 2.075 1.21 2.245 1.38 ;
      RECT 8.31 1.21 8.48 1.38 ;
      RECT 7.38 1.21 7.55 1.38 ;
      RECT 6.5 1.21 6.67 1.38 ;
      RECT 5.595 1.21 5.765 1.38 ;
      RECT 4.705 1.21 4.875 1.38 ;
      RECT 3.795 1.21 3.965 1.38 ;
      RECT 8.78 1.95 8.95 2.12 ;
      RECT 7.86 1.95 8.03 2.12 ;
      RECT 6.935 1.95 7.105 2.12 ;
      RECT 6.055 1.95 6.225 2.12 ;
      RECT 5.145 1.95 5.315 2.12 ;
      RECT 4.245 1.95 4.415 2.12 ;
      RECT 3.34 1.95 3.51 2.12 ;
      RECT 2.49 1.95 2.66 2.12 ;
      RECT 2.92 1.21 3.09 1.38 ;
      RECT 7.41 2.715 7.58 2.885 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 8.32 2.715 8.49 2.885 ;
      RECT 9.25 2.715 9.42 2.885 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.515 2.715 6.685 2.885 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.595 2.715 5.765 2.885 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.715 2.715 4.885 2.885 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.81 2.715 3.98 2.885 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.91 2.715 3.08 2.885 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.08 2.715 2.25 2.885 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
  END
END scs8ls_lpflow_clkbufkapwr_16

MACRO scs8ls_lpflow_clkbufkapwr_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.01 1.495 2.15 ;
    END
    ANTENNAGATEAREA 0.231 ;
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 0.35 0.885 0.79 ;
        RECT 0.715 0.79 0.885 1.82 ;
        RECT 0.555 1.82 0.885 2.15 ;
    END
    ANTENNADIFFAREA 0.4536 ;
  END X

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 1.85 2.945 ;
    END
  END kapwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.105 2.66 0.435 2.945 ;
      RECT 1.005 2.66 1.335 2.945 ;
      RECT 1.535 2.49 1.835 2.65 ;
      RECT 0.215 2.32 1.835 2.49 ;
      RECT 1.665 0.81 1.835 2.32 ;
      RECT 1.475 0.35 1.835 0.81 ;
      RECT 0.215 1.63 0.385 2.32 ;
      RECT 0.215 0.96 0.545 1.63 ;
      RECT 0 3.245 1.92 3.415 ;
      RECT 0 -0.085 1.92 0.085 ;
      RECT 1.055 0.085 1.305 0.81 ;
      RECT 0.115 0.085 0.365 0.79 ;
    LAYER mcon ;
      RECT 1.115 2.715 1.285 2.885 ;
      RECT 0.185 2.715 0.355 2.885 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_lpflow_clkbufkapwr_2

MACRO scs8ls_lpflow_clkbufkapwr_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.88 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.56 0.35 0.89 0.98 ;
        RECT 0.535 0.98 1.75 1.15 ;
        RECT 0.535 1.15 0.705 1.92 ;
        RECT 1.42 0.35 1.75 0.98 ;
        RECT 0.535 1.92 1.795 2.09 ;
        RECT 0.535 2.09 0.815 2.98 ;
        RECT 1.465 2.09 1.795 2.98 ;
    END
    ANTENNADIFFAREA 0.924 ;
  END X

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.055 1.08 2.455 1.41 ;
    END
    ANTENNAGATEAREA 0.231 ;
  END A

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 2.81 2.945 ;
    END
  END kapwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.88 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.88 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.995 1.92 2.245 2.98 ;
      RECT 1.015 2.26 1.295 2.98 ;
      RECT 0.115 1.82 0.365 2.98 ;
      RECT 2.415 1.75 2.795 2.98 ;
      RECT 0.875 1.58 2.795 1.75 ;
      RECT 2.625 0.81 2.795 1.58 ;
      RECT 2.42 0.48 2.795 0.81 ;
      RECT 0.875 1.35 1.885 1.58 ;
      RECT 0 3.245 2.88 3.415 ;
      RECT 0 -0.085 2.88 0.085 ;
      RECT 1.92 0.085 2.25 0.81 ;
      RECT 0.13 0.085 0.38 0.81 ;
      RECT 1.07 0.085 1.24 0.81 ;
    LAYER mcon ;
      RECT 1.115 2.715 1.285 2.885 ;
      RECT 2.075 2.715 2.245 2.885 ;
      RECT 0.155 2.715 0.325 2.885 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_lpflow_clkbufkapwr_4

MACRO scs8ls_lpflow_clkbufkapwr_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 5.28 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.095 1.78 ;
    END
    ANTENNAGATEAREA 0.462 ;
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.71 1.18 5.155 1.69 ;
        RECT 1.615 1.69 5.155 1.86 ;
        RECT 4.71 1.02 4.88 1.18 ;
        RECT 1.615 1.86 1.905 2.98 ;
        RECT 2.515 1.86 2.845 2.98 ;
        RECT 3.415 1.86 3.745 2.98 ;
        RECT 4.365 1.86 4.71 2.92 ;
        RECT 1.615 0.85 4.88 1.02 ;
        RECT 1.615 0.35 1.945 0.85 ;
        RECT 2.615 0.35 2.865 0.85 ;
        RECT 3.555 0.35 3.77 0.85 ;
        RECT 4.44 0.35 4.665 0.85 ;
    END
    ANTENNADIFFAREA 1.8417 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 5.28 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 5.28 3.575 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 5.21 2.945 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 5.28 0.085 ;
      RECT 4.835 0.085 5.165 0.68 ;
      RECT 0.115 0.085 0.445 0.81 ;
      RECT 1.115 0.085 1.445 0.81 ;
      RECT 2.115 0.085 2.445 0.68 ;
      RECT 3.045 0.085 3.375 0.68 ;
      RECT 3.94 0.085 4.27 0.68 ;
      RECT 0 3.245 5.28 3.415 ;
      RECT 4.91 2.03 5.16 2.98 ;
      RECT 3.945 2.03 4.195 2.98 ;
      RECT 3.015 2.03 3.215 2.98 ;
      RECT 2.075 2.03 2.315 2.98 ;
      RECT 1.115 2.29 1.445 2.98 ;
      RECT 0.115 1.95 0.445 2.98 ;
      RECT 1.275 1.19 4.515 1.52 ;
      RECT 0.615 2.12 0.945 2.98 ;
      RECT 0.615 1.95 1.445 2.12 ;
      RECT 1.275 1.52 1.445 1.95 ;
      RECT 1.275 1.15 1.445 1.19 ;
      RECT 0.615 0.98 1.445 1.15 ;
      RECT 0.615 0.35 0.945 0.98 ;
    LAYER mcon ;
      RECT 0.155 2.715 0.325 2.885 ;
      RECT 1.115 2.715 1.285 2.885 ;
      RECT 2.075 2.715 2.245 2.885 ;
      RECT 3.035 2.715 3.205 2.885 ;
      RECT 3.995 2.715 4.165 2.885 ;
      RECT 4.955 2.715 5.125 2.885 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_lpflow_clkbufkapwr_8

MACRO scs8ls_lpflow_clkinvkapwr_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.44 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615 0.35 1.325 0.68 ;
        RECT 1.085 0.68 1.325 2.1 ;
        RECT 0.555 2.1 1.325 2.43 ;
        RECT 0.555 2.43 0.835 3 ;
    END
    ANTENNADIFFAREA 0.47735 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.18 0.735 1.78 ;
        RECT 0.405 1.78 0.735 1.93 ;
        RECT 0.405 0.92 0.735 1.18 ;
    END
    ANTENNAGATEAREA 0.315 ;
  END A

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 1.37 2.945 ;
    END
  END kapwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.44 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.44 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.105 2.1 0.355 2.98 ;
      RECT 1.005 2.6 1.335 3.075 ;
      RECT 0 -0.085 1.44 0.085 ;
      RECT 0.115 0.085 0.445 0.75 ;
      RECT 0 3.245 1.44 3.415 ;
    LAYER mcon ;
      RECT 0.155 2.715 0.325 2.885 ;
      RECT 1.085 2.715 1.255 2.885 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_clkinvkapwr_1

MACRO scs8ls_lpflow_clkinvkapwr_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 11.52 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.01 1.18 10.48 1.41 ;
    END
    ANTENNAGATEAREA 5.04 ;
  END A

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 11.45 2.945 ;
    END
  END kapwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 11.52 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 11.52 3.575 ;
    END
  END vpwr

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.575 1.55 10.945 1.78 ;
    END
    ANTENNADIFFAREA 5.04 ;
  END Y

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER mcon ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.675 1.21 5.845 1.38 ;
      RECT 5.595 2.715 5.765 2.885 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 5.16 1.58 5.33 1.75 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.72 1.21 4.89 1.38 ;
      RECT 4.695 2.715 4.865 2.885 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 4.25 1.58 4.42 1.75 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.8 1.21 3.97 1.38 ;
      RECT 3.795 2.715 3.965 2.885 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.36 1.58 3.53 1.75 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.895 2.715 3.065 2.885 ;
      RECT 2.885 1.21 3.055 1.38 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.44 1.58 2.61 1.75 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.995 2.715 2.165 2.885 ;
      RECT 1.975 1.21 2.145 1.38 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.535 1.58 1.705 1.75 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 1.095 2.715 1.265 2.885 ;
      RECT 1.07 1.21 1.24 1.38 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 1.58 0.805 1.75 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 2.715 0.325 2.885 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 9.84 1.58 10.01 1.75 ;
      RECT 11.195 -0.085 11.365 0.085 ;
      RECT 11.195 3.245 11.365 3.415 ;
      RECT 11.155 2.715 11.325 2.885 ;
      RECT 10.715 -0.085 10.885 0.085 ;
      RECT 10.715 1.58 10.885 1.75 ;
      RECT 10.255 2.715 10.425 2.885 ;
      RECT 10.25 1.21 10.42 1.38 ;
      RECT 10.235 -0.085 10.405 0.085 ;
      RECT 10.235 3.245 10.405 3.415 ;
      RECT 9.755 -0.085 9.925 0.085 ;
      RECT 9.755 3.245 9.925 3.415 ;
      RECT 9.355 1.21 9.525 1.38 ;
      RECT 9.355 2.715 9.525 2.885 ;
      RECT 9.275 -0.085 9.445 0.085 ;
      RECT 9.275 3.245 9.445 3.415 ;
      RECT 8.92 1.58 9.09 1.75 ;
      RECT 10.715 3.245 10.885 3.415 ;
      RECT 8.795 -0.085 8.965 0.085 ;
      RECT 8.795 3.245 8.965 3.415 ;
      RECT 8.455 2.715 8.625 2.885 ;
      RECT 8.43 1.21 8.6 1.38 ;
      RECT 8.315 -0.085 8.485 0.085 ;
      RECT 8.315 3.245 8.485 3.415 ;
      RECT 8.005 1.58 8.175 1.75 ;
      RECT 7.835 -0.085 8.005 0.085 ;
      RECT 7.835 3.245 8.005 3.415 ;
      RECT 7.565 1.21 7.735 1.38 ;
      RECT 7.555 2.715 7.725 2.885 ;
      RECT 7.355 -0.085 7.525 0.085 ;
      RECT 7.355 3.245 7.525 3.415 ;
      RECT 7.095 1.58 7.265 1.75 ;
      RECT 6.875 -0.085 7.045 0.085 ;
      RECT 6.875 3.245 7.045 3.415 ;
      RECT 6.64 1.21 6.81 1.38 ;
      RECT 6.545 2.715 6.715 2.885 ;
      RECT 6.395 -0.085 6.565 0.085 ;
      RECT 6.395 3.245 6.565 3.415 ;
      RECT 6.1 1.58 6.27 1.75 ;
      RECT 5.915 -0.085 6.085 0.085 ;
    LAYER li1 ;
      RECT 6.595 1.18 6.855 1.58 ;
      RECT 6.49 1.82 6.795 2.98 ;
      RECT 9.305 1.82 9.575 2.98 ;
      RECT 6.06 1.08 6.305 2.98 ;
      RECT 6.06 0.945 6.445 1.08 ;
      RECT 6.13 0.38 6.445 0.945 ;
      RECT 9.755 1.55 10.03 2.98 ;
      RECT 5.63 1.18 5.89 1.58 ;
      RECT 5.595 1.82 5.845 2.98 ;
      RECT 5.105 1.04 5.395 2.98 ;
      RECT 5.105 0.87 5.525 1.04 ;
      RECT 5.265 0.38 5.525 0.87 ;
      RECT 4.675 1.18 4.935 1.58 ;
      RECT 4.675 1.82 4.915 2.98 ;
      RECT 4.165 1.01 4.495 2.98 ;
      RECT 4.165 0.945 4.595 1.01 ;
      RECT 4.265 0.38 4.595 0.945 ;
      RECT 10.645 1.55 10.92 2.98 ;
      RECT 3.765 1.18 3.995 1.58 ;
      RECT 11.1 1.815 11.405 2.98 ;
      RECT 7.515 1.31 7.79 1.58 ;
      RECT 7.515 1.08 10.475 1.31 ;
      RECT 8.38 1.31 8.655 1.58 ;
      RECT 9.305 1.31 9.58 1.58 ;
      RECT 10.2 1.31 10.475 1.58 ;
      RECT 8.825 1.55 9.135 2.98 ;
      RECT 8.395 1.82 8.625 2.98 ;
      RECT 7.975 1.55 8.205 2.98 ;
      RECT 7.495 1.82 7.785 2.98 ;
      RECT 7.03 0.38 7.315 2.98 ;
      RECT 3.795 1.82 3.965 2.98 ;
      RECT 3.265 0.38 3.595 2.98 ;
      RECT 2.845 1.18 3.095 1.58 ;
      RECT 2.85 1.82 3.08 2.98 ;
      RECT 0.115 0.085 0.405 0.84 ;
      RECT 0 -0.085 11.52 0.085 ;
      RECT 1.015 0.085 1.265 0.84 ;
      RECT 1.91 0.085 2.165 0.84 ;
      RECT 2.845 0.085 3.095 0.795 ;
      RECT 3.765 0.085 4.055 0.775 ;
      RECT 4.775 0.085 5.085 0.7 ;
      RECT 5.725 0.085 5.96 0.775 ;
      RECT 6.615 0.085 6.86 0.775 ;
      RECT 7.485 0.085 9.695 0.71 ;
      RECT 0 3.245 11.52 3.415 ;
      RECT 2.365 0.38 2.665 2.98 ;
      RECT 1.92 1.18 2.19 1.58 ;
      RECT 1.925 1.82 2.19 2.98 ;
      RECT 10.2 1.82 10.465 2.98 ;
      RECT 1.465 0.945 1.74 2.98 ;
      RECT 1.445 0.38 1.74 0.945 ;
      RECT 1.02 1.18 1.29 1.58 ;
      RECT 1.03 1.82 1.285 2.98 ;
      RECT 0.585 0.38 0.845 2.98 ;
      RECT 0.115 1.82 0.405 2.98 ;
  END
END scs8ls_lpflow_clkinvkapwr_16

MACRO scs8ls_lpflow_clkinvkapwr_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.35 1.315 1.78 ;
    END
    ANTENNAGATEAREA 0.63 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.18 1.795 1.95 ;
        RECT 0.12 1.95 1.795 2.12 ;
        RECT 0.615 1.01 1.795 1.18 ;
        RECT 0.12 2.12 0.45 2.98 ;
        RECT 1.02 2.12 1.35 2.98 ;
        RECT 0.615 0.51 1.305 1.01 ;
    END
    ANTENNADIFFAREA 0.994 ;
  END Y

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 1.85 2.945 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 1.55 2.29 1.8 2.98 ;
      RECT 0.62 2.29 0.82 2.98 ;
      RECT 0 3.245 1.92 3.415 ;
      RECT 0 -0.085 1.92 0.085 ;
      RECT 1.475 0.085 1.805 0.84 ;
      RECT 0.115 0.085 0.445 0.84 ;
    LAYER mcon ;
      RECT 1.595 2.715 1.765 2.885 ;
      RECT 0.635 2.715 0.805 2.885 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_lpflow_clkinvkapwr_2

MACRO scs8ls_lpflow_clkinvkapwr_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.35 2.755 1.78 ;
    END
    ANTENNAGATEAREA 1.26 ;
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.18 3.235 1.95 ;
        RECT 0.265 1.95 3.235 2.12 ;
        RECT 0.265 1.01 3.235 1.18 ;
        RECT 0.565 2.12 0.895 2.98 ;
        RECT 1.465 2.12 1.795 2.98 ;
        RECT 2.415 2.12 2.745 2.98 ;
        RECT 0.265 1.18 0.435 1.95 ;
        RECT 0.99 0.51 1.745 1.01 ;
        RECT 2.415 0.38 2.745 1.01 ;
    END
    ANTENNADIFFAREA 1.4322 ;
  END Y

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 3.29 2.945 ;
    END
  END kapwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 2.915 2.29 3.245 2.98 ;
      RECT 1.995 2.29 2.245 2.98 ;
      RECT 1.095 2.29 1.265 2.98 ;
      RECT 0.115 2.29 0.365 2.98 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.915 0.085 3.245 0.84 ;
      RECT 0.115 0.085 0.82 0.71 ;
      RECT 1.915 0.085 2.245 0.84 ;
    LAYER mcon ;
      RECT 0.155 2.715 0.325 2.885 ;
      RECT 1.095 2.715 1.265 2.885 ;
      RECT 1.995 2.715 2.165 2.885 ;
      RECT 2.995 2.715 3.165 2.885 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
  END
END scs8ls_lpflow_clkinvkapwr_4

MACRO scs8ls_lpflow_clkinvkapwr_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 6.24 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885 1.18 6.115 1.95 ;
        RECT 0.285 1.95 6.115 2.12 ;
        RECT 0.285 1.01 6.115 1.18 ;
        RECT 0.59 2.12 0.92 2.98 ;
        RECT 1.54 2.12 1.87 2.98 ;
        RECT 2.49 2.12 2.82 2.98 ;
        RECT 3.44 2.12 3.77 2.98 ;
        RECT 4.39 2.12 4.72 2.98 ;
        RECT 5.34 2.12 5.67 2.98 ;
        RECT 0.285 1.18 0.455 1.95 ;
        RECT 0.615 0.51 2.625 1.01 ;
        RECT 3.295 0.38 3.625 1.01 ;
        RECT 4.295 0.38 4.625 1.01 ;
        RECT 5.295 0.38 5.625 1.01 ;
    END
    ANTENNADIFFAREA 3.2424 ;
  END Y

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625 1.35 5.715 1.78 ;
    END
    ANTENNAGATEAREA 2.52 ;
  END A

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 6.17 2.945 ;
    END
  END kapwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 6.24 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 6.24 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.115 2.29 0.39 2.98 ;
      RECT 0 -0.085 6.24 0.085 ;
      RECT 5.795 0.085 6.125 0.84 ;
      RECT 0.115 0.085 0.445 0.84 ;
      RECT 2.795 0.085 3.125 0.84 ;
      RECT 3.795 0.085 4.125 0.84 ;
      RECT 4.795 0.085 5.125 0.84 ;
      RECT 0 3.245 6.24 3.415 ;
      RECT 5.87 2.29 6.12 2.98 ;
      RECT 4.92 2.29 5.17 2.98 ;
      RECT 3.97 2.29 4.22 2.98 ;
      RECT 3.02 2.29 3.27 2.98 ;
      RECT 2.07 2.29 2.32 2.98 ;
      RECT 1.12 2.29 1.37 2.98 ;
    LAYER mcon ;
      RECT 0.155 2.715 0.325 2.885 ;
      RECT 1.12 2.715 1.29 2.885 ;
      RECT 2.07 2.715 2.24 2.885 ;
      RECT 3.02 2.715 3.19 2.885 ;
      RECT 3.97 2.715 4.14 2.885 ;
      RECT 4.92 2.715 5.09 2.885 ;
      RECT 5.87 2.715 6.04 2.885 ;
      RECT 5.915 -0.085 6.085 0.085 ;
      RECT 5.435 -0.085 5.605 0.085 ;
      RECT 4.955 -0.085 5.125 0.085 ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 5.915 3.245 6.085 3.415 ;
      RECT 5.435 3.245 5.605 3.415 ;
      RECT 4.955 3.245 5.125 3.415 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_clkinvkapwr_8

MACRO scs8ls_lpflow_decapkapwr_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 1.92 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 1.92 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 1.92 0.245 ;
    END
  END vgnd

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 1.85 2.945 ;
    END
  END kapwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.605 0.715 0.855 1.585 ;
      RECT 0.24 0.085 0.855 0.715 ;
      RECT 0 -0.085 1.92 0.085 ;
      RECT 1.43 0.085 1.68 0.715 ;
      RECT 0 3.245 1.92 3.415 ;
      RECT 0.24 2.67 1.68 3 ;
      RECT 1.065 1.25 1.315 2.67 ;
    LAYER mcon ;
      RECT 1.21 2.725 1.38 2.895 ;
      RECT 0.85 2.725 1.02 2.895 ;
      RECT 0.49 2.725 0.66 2.895 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_decapkapwr_4

MACRO scs8ls_lpflow_decapkapwr_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.84 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN kapwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.07 2.675 3.77 2.945 ;
    END
  END kapwr

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.84 3.575 ;
    END
  END vpwr

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.84 0.245 ;
    END
  END vgnd

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.79 0.805 1.12 1.585 ;
      RECT 0.555 0.085 1.12 0.805 ;
      RECT 0 -0.085 3.84 0.085 ;
      RECT 1.755 0.085 2.085 0.805 ;
      RECT 2.66 0.085 3.28 0.805 ;
      RECT 2.66 0.805 3.065 1.58 ;
      RECT 0 3.245 3.84 3.415 ;
      RECT 0.555 2.675 3.29 2.98 ;
      RECT 0.555 2.295 0.805 2.675 ;
      RECT 3.04 2.295 3.29 2.675 ;
      RECT 1.45 1.25 2.385 2.675 ;
    LAYER mcon ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.7 2.725 2.87 2.895 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.34 2.725 2.51 2.895 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 1.98 2.725 2.15 2.895 ;
      RECT 1.62 2.725 1.79 2.895 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 3.06 2.725 3.23 2.895 ;
      RECT 1.21 2.725 1.38 2.895 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.85 2.725 1.02 2.895 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_decapkapwr_8

MACRO scs8ls_lpflow_isobufsrc_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.43 0.865 1.75 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.07 0.92 2.315 1.815 ;
        RECT 1.925 1.815 2.315 3.075 ;
        RECT 1.39 0.75 2.315 0.92 ;
        RECT 1.39 0.255 1.65 0.75 ;
    END
    ANTENNADIFFAREA 0.7075 ;
  END X

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035 1.43 1.415 1.75 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END SLEEP

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 2.4 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 2.4 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0.39 1.945 1.755 2.14 ;
      RECT 1.585 1.55 1.755 1.945 ;
      RECT 1.585 1.26 1.9 1.55 ;
      RECT 0.355 1.09 1.9 1.26 ;
      RECT 0.355 0.35 0.625 1.09 ;
      RECT 0 -0.085 2.4 0.085 ;
      RECT 1.82 0.085 2.15 0.58 ;
      RECT 0.795 0.085 1.125 0.58 ;
      RECT 0 3.245 2.4 3.415 ;
      RECT 0.96 2.31 1.29 3.245 ;
    LAYER mcon ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_isobufsrc_1

MACRO scs8ls_lpflow_isobufsrc_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 3.36 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055 1.26 1.775 1.47 ;
        RECT 1.055 1.09 2.805 1.26 ;
        RECT 2.555 1.26 2.805 1.55 ;
    END
    ANTENNAGATEAREA 0.558 ;
  END SLEEP

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555 1.21 0.885 1.515 ;
    END
    ANTENNAGATEAREA 0.126 ;
  END A

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.015 0.92 3.275 1.72 ;
        RECT 2.445 1.72 3.275 1.95 ;
        RECT 1.435 0.75 3.275 0.92 ;
        RECT 2.445 1.95 2.615 2.025 ;
        RECT 1.435 0.58 1.695 0.75 ;
        RECT 2.365 0.58 2.555 0.75 ;
        RECT 1.82 2.025 2.615 2.195 ;
        RECT 1.82 2.195 2.07 2.725 ;
    END
    ANTENNADIFFAREA 0.7504 ;
  END X

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 3.36 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 3.36 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 -0.085 3.36 0.085 ;
      RECT 2.725 0.085 3.055 0.58 ;
      RECT 0.59 0.97 0.895 1.015 ;
      RECT 0.59 0.94 0.93 0.97 ;
      RECT 0.59 0.885 0.965 0.94 ;
      RECT 0.59 0.085 1.265 0.885 ;
      RECT 1.865 0.085 2.195 0.58 ;
      RECT 0.16 1.685 2.275 1.855 ;
      RECT 1.945 1.43 2.275 1.685 ;
      RECT 0.16 1.855 0.6 2.21 ;
      RECT 0.16 1.03 0.385 1.685 ;
      RECT 0.16 0.7 0.41 1.03 ;
      RECT 1.395 2.895 2.6 3.075 ;
      RECT 2.27 2.365 2.6 2.895 ;
      RECT 1.395 2.025 1.625 2.895 ;
      RECT 0 3.245 3.36 3.415 ;
      RECT 2.79 2.3 3.05 3.245 ;
      RECT 0.875 2.025 1.225 3.245 ;
    LAYER mcon ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_isobufsrc_2

MACRO scs8ls_lpflow_isobufsrc_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 3.33 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.475 0.92 4.7 2.035 ;
        RECT 1.615 2.035 4.7 2.205 ;
        RECT 1.2 0.75 4.7 0.92 ;
        RECT 1.615 2.205 1.945 2.235 ;
        RECT 3.415 2.205 3.745 2.58 ;
        RECT 1.2 0.645 1.46 0.75 ;
        RECT 2.13 0.645 2.32 0.75 ;
        RECT 2.99 0.625 3.18 0.75 ;
        RECT 3.86 0.625 4.03 0.75 ;
    END
    ANTENNADIFFAREA 1.5156 ;
  END X

  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.065 1.43 2.725 1.695 ;
        RECT 0.925 1.695 4.305 1.865 ;
        RECT 0.925 1.43 1.255 1.695 ;
        RECT 4.045 1.22 4.305 1.695 ;
    END
    ANTENNAGATEAREA 1.116 ;
  END SLEEP

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.345 0.415 1.76 ;
    END
    ANTENNAGATEAREA 0.279 ;
  END A

  PIN vgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 -0.245 4.8 0.245 ;
    END
  END vgnd

  PIN vpwr
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 3.085 4.8 3.575 ;
    END
  END vpwr

  PIN vpb
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0 3.08 0.25 3.33 ;
    END
  END vpb

  PIN vnb
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0 0 0.25 0.25 ;
    END
  END vnb
  OBS
    LAYER li1 ;
      RECT 0 3.245 4.8 3.415 ;
      RECT 4.315 2.375 4.645 3.245 ;
      RECT 2.515 2.745 2.845 3.245 ;
      RECT 0.555 2.27 0.835 3.245 ;
      RECT 0 -0.085 4.8 0.085 ;
      RECT 4.23 0.085 4.56 0.58 ;
      RECT 0.69 0.085 1.02 0.835 ;
      RECT 1.63 0.085 1.96 0.58 ;
      RECT 2.49 0.085 2.82 0.58 ;
      RECT 3.35 0.085 3.68 0.58 ;
      RECT 3.045 2.75 4.125 2.92 ;
      RECT 3.935 2.375 4.125 2.75 ;
      RECT 1.075 2.575 1.325 3 ;
      RECT 1.075 2.035 1.335 2.405 ;
      RECT 1.075 2.405 3.215 2.575 ;
      RECT 2.145 2.575 2.315 2.995 ;
      RECT 3.045 2.575 3.215 2.75 ;
      RECT 3.045 2.375 3.215 2.405 ;
      RECT 0.585 1.175 3.635 1.26 ;
      RECT 3.305 1.26 3.635 1.515 ;
      RECT 0.26 1.09 3.635 1.175 ;
      RECT 0.1 2.1 0.37 3.075 ;
      RECT 0.1 1.93 0.755 2.1 ;
      RECT 0.585 1.26 0.755 1.93 ;
      RECT 0.26 1.005 0.785 1.09 ;
      RECT 0.26 0.255 0.52 1.005 ;
      RECT 1.565 1.26 1.895 1.515 ;
    LAYER mcon ;
      RECT 4.475 -0.085 4.645 0.085 ;
      RECT 4.475 3.245 4.645 3.415 ;
      RECT 3.995 -0.085 4.165 0.085 ;
      RECT 3.995 3.245 4.165 3.415 ;
      RECT 3.515 -0.085 3.685 0.085 ;
      RECT 3.515 3.245 3.685 3.415 ;
      RECT 3.035 -0.085 3.205 0.085 ;
      RECT 3.035 3.245 3.205 3.415 ;
      RECT 2.555 -0.085 2.725 0.085 ;
      RECT 2.555 3.245 2.725 3.415 ;
      RECT 2.075 -0.085 2.245 0.085 ;
      RECT 2.075 3.245 2.245 3.415 ;
      RECT 1.595 -0.085 1.765 0.085 ;
      RECT 1.595 3.245 1.765 3.415 ;
      RECT 1.115 -0.085 1.285 0.085 ;
      RECT 1.115 3.245 1.285 3.415 ;
      RECT 0.635 -0.085 0.805 0.085 ;
      RECT 0.635 3.245 0.805 3.415 ;
      RECT 0.155 -0.085 0.325 0.085 ;
      RECT 0.155 3.245 0.325 3.415 ;
  END
END scs8ls_lpflow_isobufsrc_4
  
END LIBRARY
